* EQUIVALENT CIRCUIT FOR VECTOR FITTED
* Created by wyz
*
.SUBCKT s_equivalent p1 p2
*
* Port network for port 1
V1 p1 s1 0
R1 s1 0 50.0
Gd1_1 0 s1 p1 0 -0.019262662535517755
Fd1_1 0 s1 V1 -0.9631331267758878
Gr1_1_1 0 s1 x1_a1 0 -22512084776.36006
Gr2_re_1_1 0 s1 x2_re_a1 0 20420362323.016293
Gr2_im_1_1 0 s1 x2_im_a1 0 2972214744.9561706
Gd1_2 0 s1 p2 0 -0.0016343936673183504
Fd1_2 0 s1 V2 -0.08171968336591752
Gr1_1_2 0 s1 x1_a2 0 8983926499.253344
Gr2_re_1_2 0 s1 x2_re_a2 0 22937049642.695232
Gr2_im_1_2 0 s1 x2_im_a2 0 -1691112963.819676
*
* State networks driven by port 1
Cx1_a1 x1_a1 0 1.0
Gx1_a1 0 x1_a1 p1 0 0.07071067811865475
Fx1_a1 0 x1_a1 V1 3.5355339059327378
Rp1_a1 0 x1_a1 4.439606360475265e-13
Cx2_re_a1 x2_re_a1 0 1.0
Gx2_re_a1 0 x2_re_a1 p1 0 0.1414213562373095
Fx2_re_a1 0 x2_re_a1 V1 7.0710678118654755
Rp2_re_re_a1 0 x2_re_a1 1.2563049453689557e-11
Gp2_re_im_a1 0 x2_re_a1 x2_im_a1 0 533476609939.1895
Cx2_im_a1 x2_im_a1 0 1.0
Gp2_im_re_a1 0 x2_im_a1 x2_re_a1 0 -533476609939.1895
Rp2_im_im_a1 0 x2_im_a1 1.2563049453689557e-11
*
* Port network for port 2
V2 p2 s2 0
R2 s2 0 50.0
Gd2_1 0 s2 p1 0 -0.0016343940302883653
Fd2_1 0 s2 V1 -0.08171970151441828
Gr1_2_1 0 s2 x1_a1 0 8983926498.965857
Gr2_re_2_1 0 s2 x2_re_a1 0 22937049669.817776
Gr2_im_2_1 0 s2 x2_im_a1 0 -1691113010.291936
Gd2_2 0 s2 p2 0 0.0187133623188902
Fd2_2 0 s2 V2 0.93566811594451
Gr1_2_2 0 s2 x1_a2 0 -1324757794605.9355
Gr2_re_2_2 0 s2 x2_re_a2 0 24287089530.553734
Gr2_im_2_2 0 s2 x2_im_a2 0 -7538139793.597747
*
* State networks driven by port 2
Cx1_a2 x1_a2 0 1.0
Gx1_a2 0 x1_a2 p2 0 0.07071067811865475
Fx1_a2 0 x1_a2 V2 3.5355339059327378
Rp1_a2 0 x1_a2 4.439606360475265e-13
Cx2_re_a2 x2_re_a2 0 1.0
Gx2_re_a2 0 x2_re_a2 p2 0 0.1414213562373095
Fx2_re_a2 0 x2_re_a2 V2 7.0710678118654755
Rp2_re_re_a2 0 x2_re_a2 1.2563049453689557e-11
Gp2_re_im_a2 0 x2_re_a2 x2_im_a2 0 533476609939.1895
Cx2_im_a2 x2_im_a2 0 1.0
Gp2_im_re_a2 0 x2_im_a2 x2_re_a2 0 -533476609939.1895
Rp2_im_im_a2 0 x2_im_a2 1.2563049453689557e-11
.ENDS s_equivalent
