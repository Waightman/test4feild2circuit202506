* EQUIVALENT CIRCUIT FOR VECTOR FITTED
* Created by wyz
*
.SUBCKT s_equivalent p1 p2
*
* Port network for port 1
V1 p1 s1 0
R1 s1 0 50.0
Gd1_1 0 s1 p1 0 0.0003110693704729122
Fd1_1 0 s1 V1 0.01555346852364561
Gr1_1_1 0 s1 x1_a1 0 -3368187027.594035
Gr2_re_1_1 0 s1 x2_re_a1 0 -30766869.066676043
Gr2_im_1_1 0 s1 x2_im_a1 0 100392901.51010174
Gr3_re_1_1 0 s1 x3_re_a1 0 3262428537.608702
Gr3_im_1_1 0 s1 x3_im_a1 0 4638282076.006712
Gr4_re_1_1 0 s1 x4_re_a1 0 -4399897721.094303
Gr4_im_1_1 0 s1 x4_im_a1 0 -8136353477.688546
Gr5_re_1_1 0 s1 x5_re_a1 0 194887.43443422127
Gr5_im_1_1 0 s1 x5_im_a1 0 30614.601410188465
Gr6_re_1_1 0 s1 x6_re_a1 0 168054.8042040786
Gr6_im_1_1 0 s1 x6_im_a1 0 208186.61452473744
Gr7_re_1_1 0 s1 x7_re_a1 0 -142376467.8772501
Gr7_im_1_1 0 s1 x7_im_a1 0 -1778734115.6796474
Gr8_re_1_1 0 s1 x8_re_a1 0 900712532.6898531
Gr8_im_1_1 0 s1 x8_im_a1 0 266188716.32368398
Gr9_re_1_1 0 s1 x9_re_a1 0 -382864080.64300835
Gr9_im_1_1 0 s1 x9_im_a1 0 296593399.290862
Gr10_re_1_1 0 s1 x10_re_a1 0 2317861.5012086863
Gr10_im_1_1 0 s1 x10_im_a1 0 -3423674.5108741857
Gr11_re_1_1 0 s1 x11_re_a1 0 -314495.9788154342
Gr11_im_1_1 0 s1 x11_im_a1 0 -1308584.673824057
Gr12_re_1_1 0 s1 x12_re_a1 0 270816281.0595158
Gr12_im_1_1 0 s1 x12_im_a1 0 -803431878.679809
Gr13_re_1_1 0 s1 x13_re_a1 0 383906249.46809435
Gr13_im_1_1 0 s1 x13_im_a1 0 754515974.4450386
Gr14_re_1_1 0 s1 x14_re_a1 0 213088295.5059075
Gr14_im_1_1 0 s1 x14_im_a1 0 -592654662.4520757
Gr15_re_1_1 0 s1 x15_re_a1 0 1962934250.172265
Gr15_im_1_1 0 s1 x15_im_a1 0 1954346430.0687664
Gr16_re_1_1 0 s1 x16_re_a1 0 880187.777989353
Gr16_im_1_1 0 s1 x16_im_a1 0 -76246184.8403165
Gr17_re_1_1 0 s1 x17_re_a1 0 199737789.85648456
Gr17_im_1_1 0 s1 x17_im_a1 0 -852593629.4591384
Gd1_2 0 s1 p2 0 0.0008880606688733853
Fd1_2 0 s1 V2 0.04440303344366926
Gr1_1_2 0 s1 x1_a2 0 -10402598898.868498
Gr2_re_1_2 0 s1 x2_re_a2 0 -736374544.752954
Gr2_im_1_2 0 s1 x2_im_a2 0 -772196657.9494315
Gr3_re_1_2 0 s1 x3_re_a2 0 319920922.13839763
Gr3_im_1_2 0 s1 x3_im_a2 0 185491484.38332742
Gr4_re_1_2 0 s1 x4_re_a2 0 44561211.03510773
Gr4_im_1_2 0 s1 x4_im_a2 0 -795840506.9496604
Gr5_re_1_2 0 s1 x5_re_a2 0 -8557431.57335654
Gr5_im_1_2 0 s1 x5_im_a2 0 15614054.798876971
Gr6_re_1_2 0 s1 x6_re_a2 0 -9736471.028745988
Gr6_im_1_2 0 s1 x6_im_a2 0 1202644.3076369695
Gr7_re_1_2 0 s1 x7_re_a2 0 446218689.3404745
Gr7_im_1_2 0 s1 x7_im_a2 0 371562708.8664752
Gr8_re_1_2 0 s1 x8_re_a2 0 -2948522305.295996
Gr8_im_1_2 0 s1 x8_im_a2 0 1851155065.5306096
Gr9_re_1_2 0 s1 x9_re_a2 0 76191097.70774908
Gr9_im_1_2 0 s1 x9_im_a2 0 50848005.13096265
Gr10_re_1_2 0 s1 x10_re_a2 0 -335765.90712474234
Gr10_im_1_2 0 s1 x10_im_a2 0 -154577.25647844438
Gr11_re_1_2 0 s1 x11_re_a2 0 8147747.79816226
Gr11_im_1_2 0 s1 x11_im_a2 0 -22992198.453187883
Gr12_re_1_2 0 s1 x12_re_a2 0 6348260477.279809
Gr12_im_1_2 0 s1 x12_im_a2 0 -1590104490.5462964
Gr13_re_1_2 0 s1 x13_re_a2 0 -177535352.8464971
Gr13_im_1_2 0 s1 x13_im_a2 0 137358499.56066585
Gr14_re_1_2 0 s1 x14_re_a2 0 -3123494938.22666
Gr14_im_1_2 0 s1 x14_im_a2 0 13431169.122418571
Gr15_re_1_2 0 s1 x15_re_a2 0 158488666.80550125
Gr15_im_1_2 0 s1 x15_im_a2 0 685717696.6429961
Gr16_re_1_2 0 s1 x16_re_a2 0 318203012.5075078
Gr16_im_1_2 0 s1 x16_im_a2 0 -507208510.6569406
Gr17_re_1_2 0 s1 x17_re_a2 0 143393963.75206065
Gr17_im_1_2 0 s1 x17_im_a2 0 -116731155.66132578
*
* State networks driven by port 1
Cx1_a1 x1_a1 0 1.0
Gx1_a1 0 x1_a1 p1 0 0.07071067811865475
Fx1_a1 0 x1_a1 V1 3.5355339059327378
Rp1_a1 0 x1_a1 3.320472266722773e-12
Cx2_re_a1 x2_re_a1 0 1.0
Gx2_re_a1 0 x2_re_a1 p1 0 0.1414213562373095
Fx2_re_a1 0 x2_re_a1 V1 7.0710678118654755
Rp2_re_re_a1 0 x2_re_a1 1.222628454118507e-10
Gp2_re_im_a1 0 x2_re_a1 x2_im_a1 0 206564125909.31366
Cx2_im_a1 x2_im_a1 0 1.0
Gp2_im_re_a1 0 x2_im_a1 x2_re_a1 0 -206564125909.31366
Rp2_im_im_a1 0 x2_im_a1 1.222628454118507e-10
Cx3_re_a1 x3_re_a1 0 1.0
Gx3_re_a1 0 x3_re_a1 p1 0 0.1414213562373095
Fx3_re_a1 0 x3_re_a1 V1 7.0710678118654755
Rp3_re_re_a1 0 x3_re_a1 7.026662594154148e-11
Gp3_re_im_a1 0 x3_re_a1 x3_im_a1 0 194277309617.66318
Cx3_im_a1 x3_im_a1 0 1.0
Gp3_im_re_a1 0 x3_im_a1 x3_re_a1 0 -194277309617.66318
Rp3_im_im_a1 0 x3_im_a1 7.026662594154148e-11
Cx4_re_a1 x4_re_a1 0 1.0
Gx4_re_a1 0 x4_re_a1 p1 0 0.1414213562373095
Fx4_re_a1 0 x4_re_a1 V1 7.0710678118654755
Rp4_re_re_a1 0 x4_re_a1 4.34339120967275e-11
Gp4_re_im_a1 0 x4_re_a1 x4_im_a1 0 127783819533.63753
Cx4_im_a1 x4_im_a1 0 1.0
Gp4_im_re_a1 0 x4_im_a1 x4_re_a1 0 -127783819533.63753
Rp4_im_im_a1 0 x4_im_a1 4.34339120967275e-11
Cx5_re_a1 x5_re_a1 0 1.0
Gx5_re_a1 0 x5_re_a1 p1 0 0.1414213562373095
Fx5_re_a1 0 x5_re_a1 V1 7.0710678118654755
Rp5_re_re_a1 0 x5_re_a1 3.9241855220809974e-10
Gp5_re_im_a1 0 x5_re_a1 x5_im_a1 0 183851444273.21875
Cx5_im_a1 x5_im_a1 0 1.0
Gp5_im_re_a1 0 x5_im_a1 x5_re_a1 0 -183851444273.21875
Rp5_im_im_a1 0 x5_im_a1 3.9241855220809974e-10
Cx6_re_a1 x6_re_a1 0 1.0
Gx6_re_a1 0 x6_re_a1 p1 0 0.1414213562373095
Fx6_re_a1 0 x6_re_a1 V1 7.0710678118654755
Rp6_re_re_a1 0 x6_re_a1 5.732214204378206e-10
Gp6_re_im_a1 0 x6_re_a1 x6_im_a1 0 130040083838.637
Cx6_im_a1 x6_im_a1 0 1.0
Gp6_im_re_a1 0 x6_im_a1 x6_re_a1 0 -130040083838.637
Rp6_im_im_a1 0 x6_im_a1 5.732214204378206e-10
Cx7_re_a1 x7_re_a1 0 1.0
Gx7_re_a1 0 x7_re_a1 p1 0 0.1414213562373095
Fx7_re_a1 0 x7_re_a1 V1 7.0710678118654755
Rp7_re_re_a1 0 x7_re_a1 1.6234265289688375e-10
Gp7_re_im_a1 0 x7_re_a1 x7_im_a1 0 176597803098.30023
Cx7_im_a1 x7_im_a1 0 1.0
Gp7_im_re_a1 0 x7_im_a1 x7_re_a1 0 -176597803098.30023
Rp7_im_im_a1 0 x7_im_a1 1.6234265289688375e-10
Cx8_re_a1 x8_re_a1 0 1.0
Gx8_re_a1 0 x8_re_a1 p1 0 0.1414213562373095
Fx8_re_a1 0 x8_re_a1 V1 7.0710678118654755
Rp8_re_re_a1 0 x8_re_a1 1.4083143320865588e-10
Gp8_re_im_a1 0 x8_re_a1 x8_im_a1 0 175562128496.72046
Cx8_im_a1 x8_im_a1 0 1.0
Gp8_im_re_a1 0 x8_im_a1 x8_re_a1 0 -175562128496.72046
Rp8_im_im_a1 0 x8_im_a1 1.4083143320865588e-10
Cx9_re_a1 x9_re_a1 0 1.0
Gx9_re_a1 0 x9_re_a1 p1 0 0.1414213562373095
Fx9_re_a1 0 x9_re_a1 V1 7.0710678118654755
Rp9_re_re_a1 0 x9_re_a1 1.715215055825635e-10
Gp9_re_im_a1 0 x9_re_a1 x9_im_a1 0 170388268279.49786
Cx9_im_a1 x9_im_a1 0 1.0
Gp9_im_re_a1 0 x9_im_a1 x9_re_a1 0 -170388268279.49786
Rp9_im_im_a1 0 x9_im_a1 1.715215055825635e-10
Cx10_re_a1 x10_re_a1 0 1.0
Gx10_re_a1 0 x10_re_a1 p1 0 0.1414213562373095
Fx10_re_a1 0 x10_re_a1 V1 7.0710678118654755
Rp10_re_re_a1 0 x10_re_a1 1.279330633293622e-09
Gp10_re_im_a1 0 x10_re_a1 x10_im_a1 0 138925213075.38348
Cx10_im_a1 x10_im_a1 0 1.0
Gp10_im_re_a1 0 x10_im_a1 x10_re_a1 0 -138925213075.38348
Rp10_im_im_a1 0 x10_im_a1 1.279330633293622e-09
Cx11_re_a1 x11_re_a1 0 1.0
Gx11_re_a1 0 x11_re_a1 p1 0 0.1414213562373095
Fx11_re_a1 0 x11_re_a1 V1 7.0710678118654755
Rp11_re_re_a1 0 x11_re_a1 3.9059155840864643e-10
Gp11_re_im_a1 0 x11_re_a1 x11_im_a1 0 139719166370.31833
Cx11_im_a1 x11_im_a1 0 1.0
Gp11_im_re_a1 0 x11_im_a1 x11_re_a1 0 -139719166370.31833
Rp11_im_im_a1 0 x11_im_a1 3.9059155840864643e-10
Cx12_re_a1 x12_re_a1 0 1.0
Gx12_re_a1 0 x12_re_a1 p1 0 0.1414213562373095
Fx12_re_a1 0 x12_re_a1 V1 7.0710678118654755
Rp12_re_re_a1 0 x12_re_a1 1.049749481959773e-10
Gp12_re_im_a1 0 x12_re_a1 x12_im_a1 0 162806930635.2914
Cx12_im_a1 x12_im_a1 0 1.0
Gp12_im_re_a1 0 x12_im_a1 x12_re_a1 0 -162806930635.2914
Rp12_im_im_a1 0 x12_im_a1 1.049749481959773e-10
Cx13_re_a1 x13_re_a1 0 1.0
Gx13_re_a1 0 x13_re_a1 p1 0 0.1414213562373095
Fx13_re_a1 0 x13_re_a1 V1 7.0710678118654755
Rp13_re_re_a1 0 x13_re_a1 1.731638893406368e-10
Gp13_re_im_a1 0 x13_re_a1 x13_im_a1 0 161735038737.64923
Cx13_im_a1 x13_im_a1 0 1.0
Gp13_im_re_a1 0 x13_im_a1 x13_re_a1 0 -161735038737.64923
Rp13_im_im_a1 0 x13_im_a1 1.731638893406368e-10
Cx14_re_a1 x14_re_a1 0 1.0
Gx14_re_a1 0 x14_re_a1 p1 0 0.1414213562373095
Fx14_re_a1 0 x14_re_a1 V1 7.0710678118654755
Rp14_re_re_a1 0 x14_re_a1 1.5904302621228683e-10
Gp14_re_im_a1 0 x14_re_a1 x14_im_a1 0 154094455422.17636
Cx14_im_a1 x14_im_a1 0 1.0
Gp14_im_re_a1 0 x14_im_a1 x14_re_a1 0 -154094455422.17636
Rp14_im_im_a1 0 x14_im_a1 1.5904302621228683e-10
Cx15_re_a1 x15_re_a1 0 1.0
Gx15_re_a1 0 x15_re_a1 p1 0 0.1414213562373095
Fx15_re_a1 0 x15_re_a1 V1 7.0710678118654755
Rp15_re_re_a1 0 x15_re_a1 1.5963175233460748e-10
Gp15_re_im_a1 0 x15_re_a1 x15_im_a1 0 151958412904.65485
Cx15_im_a1 x15_im_a1 0 1.0
Gp15_im_re_a1 0 x15_im_a1 x15_re_a1 0 -151958412904.65485
Rp15_im_im_a1 0 x15_im_a1 1.5963175233460748e-10
Cx16_re_a1 x16_re_a1 0 1.0
Gx16_re_a1 0 x16_re_a1 p1 0 0.1414213562373095
Fx16_re_a1 0 x16_re_a1 V1 7.0710678118654755
Rp16_re_re_a1 0 x16_re_a1 4.085517959442536e-10
Gp16_re_im_a1 0 x16_re_a1 x16_im_a1 0 150304807574.39594
Cx16_im_a1 x16_im_a1 0 1.0
Gp16_im_re_a1 0 x16_im_a1 x16_re_a1 0 -150304807574.39594
Rp16_im_im_a1 0 x16_im_a1 4.085517959442536e-10
Cx17_re_a1 x17_re_a1 0 1.0
Gx17_re_a1 0 x17_re_a1 p1 0 0.1414213562373095
Fx17_re_a1 0 x17_re_a1 V1 7.0710678118654755
Rp17_re_re_a1 0 x17_re_a1 3.8552133160375805e-10
Gp17_re_im_a1 0 x17_re_a1 x17_im_a1 0 150713612315.05786
Cx17_im_a1 x17_im_a1 0 1.0
Gp17_im_re_a1 0 x17_im_a1 x17_re_a1 0 -150713612315.05786
Rp17_im_im_a1 0 x17_im_a1 3.8552133160375805e-10
*
* Port network for port 2
V2 p2 s2 0
R2 s2 0 50.0
Gd2_1 0 s2 p1 0 0.0008880606688730646
Fd2_1 0 s2 V1 0.044403033443653234
Gr1_2_1 0 s2 x1_a1 0 -10402598898.863747
Gr2_re_2_1 0 s2 x2_re_a1 0 -736374544.7531635
Gr2_im_2_1 0 s2 x2_im_a1 0 -772196657.9495612
Gr3_re_2_1 0 s2 x3_re_a1 0 319920922.13817346
Gr3_im_2_1 0 s2 x3_im_a1 0 185491484.38355702
Gr4_re_2_1 0 s2 x4_re_a1 0 44561211.035196215
Gr4_im_2_1 0 s2 x4_im_a1 0 -795840506.9494897
Gr5_re_2_1 0 s2 x5_re_a1 0 -8557431.573358634
Gr5_im_2_1 0 s2 x5_im_a1 0 15614054.798876785
Gr6_re_2_1 0 s2 x6_re_a1 0 -9736471.028745329
Gr6_im_2_1 0 s2 x6_im_a1 0 1202644.307636511
Gr7_re_2_1 0 s2 x7_re_a1 0 446218689.3405445
Gr7_im_2_1 0 s2 x7_im_a1 0 371562708.86629975
Gr8_re_2_1 0 s2 x8_re_a1 0 -2948522305.296232
Gr8_im_2_1 0 s2 x8_im_a1 0 1851155065.5308654
Gr9_re_2_1 0 s2 x9_re_a1 0 76191097.70776573
Gr9_im_2_1 0 s2 x9_im_a1 0 50848005.13101999
Gr10_re_2_1 0 s2 x10_re_a1 0 -335765.9071252678
Gr10_im_2_1 0 s2 x10_im_a1 0 -154577.25647877657
Gr11_re_2_1 0 s2 x11_re_a1 0 8147747.798163875
Gr11_im_2_1 0 s2 x11_im_a1 0 -22992198.453186795
Gr12_re_2_1 0 s2 x12_re_a1 0 6348260477.279915
Gr12_im_2_1 0 s2 x12_im_a1 0 -1590104490.5460944
Gr13_re_2_1 0 s2 x13_re_a1 0 -177535352.8465156
Gr13_im_2_1 0 s2 x13_im_a1 0 137358499.56062448
Gr14_re_2_1 0 s2 x14_re_a1 0 -3123494938.2267656
Gr14_im_2_1 0 s2 x14_im_a1 0 13431169.122443844
Gr15_re_2_1 0 s2 x15_re_a1 0 158488666.80568242
Gr15_im_2_1 0 s2 x15_im_a1 0 685717696.6430213
Gr16_re_2_1 0 s2 x16_re_a1 0 318203012.5075046
Gr16_im_2_1 0 s2 x16_im_a1 0 -507208510.65688425
Gr17_re_2_1 0 s2 x17_re_a1 0 143393963.75203305
Gr17_im_2_1 0 s2 x17_im_a1 0 -116731155.66138902
Gd2_2 0 s2 p2 0 0.00033354056051843923
Fd2_2 0 s2 V2 0.016677028025921962
Gr1_2_2 0 s2 x1_a2 0 -2998907055.678349
Gr2_re_2_2 0 s2 x2_re_a2 0 -12927240.519722272
Gr2_im_2_2 0 s2 x2_im_a2 0 79467423.38936985
Gr3_re_2_2 0 s2 x3_re_a2 0 3211001844.7735095
Gr3_im_2_2 0 s2 x3_im_a2 0 4595596667.802097
Gr4_re_2_2 0 s2 x4_re_a2 0 -4335935860.012611
Gr4_im_2_2 0 s2 x4_im_a2 0 -8098139912.8550005
Gr5_re_2_2 0 s2 x5_re_a2 0 -111680.77464141163
Gr5_im_2_2 0 s2 x5_im_a2 0 157089.69332840497
Gr6_re_2_2 0 s2 x6_re_a2 0 -348825.7115814165
Gr6_im_2_2 0 s2 x6_im_a2 0 -294190.30402653833
Gr7_re_2_2 0 s2 x7_re_a2 0 -98806737.48264237
Gr7_im_2_2 0 s2 x7_im_a2 0 -1773120864.8938992
Gr8_re_2_2 0 s2 x8_re_a2 0 834763680.7297922
Gr8_im_2_2 0 s2 x8_im_a2 0 215079972.47193143
Gr9_re_2_2 0 s2 x9_re_a2 0 -401237370.9491654
Gr9_im_2_2 0 s2 x9_im_a2 0 299554979.58290166
Gr10_re_2_2 0 s2 x10_re_a2 0 2148514.9239008212
Gr10_im_2_2 0 s2 x10_im_a2 0 -3581354.9523958676
Gr11_re_2_2 0 s2 x11_re_a2 0 -7147.429289976264
Gr11_im_2_2 0 s2 x11_im_a2 0 733991.6056657406
Gr12_re_2_2 0 s2 x12_re_a2 0 126021110.1311365
Gr12_im_2_2 0 s2 x12_im_a2 0 -777200505.6826302
Gr13_re_2_2 0 s2 x13_re_a2 0 410056204.91540384
Gr13_im_2_2 0 s2 x13_im_a2 0 769687399.5843744
Gr14_re_2_2 0 s2 x14_re_a2 0 103751417.42875153
Gr14_im_2_2 0 s2 x14_im_a2 0 -503610765.42559785
Gr15_re_2_2 0 s2 x15_re_a2 0 2128824834.025204
Gr15_im_2_2 0 s2 x15_im_a2 0 1934460320.568906
Gr16_re_2_2 0 s2 x16_re_a2 0 19007471.738271806
Gr16_im_2_2 0 s2 x16_im_a2 0 -45037697.957206614
Gr17_re_2_2 0 s2 x17_re_a2 0 163670435.87085682
Gr17_im_2_2 0 s2 x17_im_a2 0 -871709689.5693338
*
* State networks driven by port 2
Cx1_a2 x1_a2 0 1.0
Gx1_a2 0 x1_a2 p2 0 0.07071067811865475
Fx1_a2 0 x1_a2 V2 3.5355339059327378
Rp1_a2 0 x1_a2 3.320472266722773e-12
Cx2_re_a2 x2_re_a2 0 1.0
Gx2_re_a2 0 x2_re_a2 p2 0 0.1414213562373095
Fx2_re_a2 0 x2_re_a2 V2 7.0710678118654755
Rp2_re_re_a2 0 x2_re_a2 1.222628454118507e-10
Gp2_re_im_a2 0 x2_re_a2 x2_im_a2 0 206564125909.31366
Cx2_im_a2 x2_im_a2 0 1.0
Gp2_im_re_a2 0 x2_im_a2 x2_re_a2 0 -206564125909.31366
Rp2_im_im_a2 0 x2_im_a2 1.222628454118507e-10
Cx3_re_a2 x3_re_a2 0 1.0
Gx3_re_a2 0 x3_re_a2 p2 0 0.1414213562373095
Fx3_re_a2 0 x3_re_a2 V2 7.0710678118654755
Rp3_re_re_a2 0 x3_re_a2 7.026662594154148e-11
Gp3_re_im_a2 0 x3_re_a2 x3_im_a2 0 194277309617.66318
Cx3_im_a2 x3_im_a2 0 1.0
Gp3_im_re_a2 0 x3_im_a2 x3_re_a2 0 -194277309617.66318
Rp3_im_im_a2 0 x3_im_a2 7.026662594154148e-11
Cx4_re_a2 x4_re_a2 0 1.0
Gx4_re_a2 0 x4_re_a2 p2 0 0.1414213562373095
Fx4_re_a2 0 x4_re_a2 V2 7.0710678118654755
Rp4_re_re_a2 0 x4_re_a2 4.34339120967275e-11
Gp4_re_im_a2 0 x4_re_a2 x4_im_a2 0 127783819533.63753
Cx4_im_a2 x4_im_a2 0 1.0
Gp4_im_re_a2 0 x4_im_a2 x4_re_a2 0 -127783819533.63753
Rp4_im_im_a2 0 x4_im_a2 4.34339120967275e-11
Cx5_re_a2 x5_re_a2 0 1.0
Gx5_re_a2 0 x5_re_a2 p2 0 0.1414213562373095
Fx5_re_a2 0 x5_re_a2 V2 7.0710678118654755
Rp5_re_re_a2 0 x5_re_a2 3.9241855220809974e-10
Gp5_re_im_a2 0 x5_re_a2 x5_im_a2 0 183851444273.21875
Cx5_im_a2 x5_im_a2 0 1.0
Gp5_im_re_a2 0 x5_im_a2 x5_re_a2 0 -183851444273.21875
Rp5_im_im_a2 0 x5_im_a2 3.9241855220809974e-10
Cx6_re_a2 x6_re_a2 0 1.0
Gx6_re_a2 0 x6_re_a2 p2 0 0.1414213562373095
Fx6_re_a2 0 x6_re_a2 V2 7.0710678118654755
Rp6_re_re_a2 0 x6_re_a2 5.732214204378206e-10
Gp6_re_im_a2 0 x6_re_a2 x6_im_a2 0 130040083838.637
Cx6_im_a2 x6_im_a2 0 1.0
Gp6_im_re_a2 0 x6_im_a2 x6_re_a2 0 -130040083838.637
Rp6_im_im_a2 0 x6_im_a2 5.732214204378206e-10
Cx7_re_a2 x7_re_a2 0 1.0
Gx7_re_a2 0 x7_re_a2 p2 0 0.1414213562373095
Fx7_re_a2 0 x7_re_a2 V2 7.0710678118654755
Rp7_re_re_a2 0 x7_re_a2 1.6234265289688375e-10
Gp7_re_im_a2 0 x7_re_a2 x7_im_a2 0 176597803098.30023
Cx7_im_a2 x7_im_a2 0 1.0
Gp7_im_re_a2 0 x7_im_a2 x7_re_a2 0 -176597803098.30023
Rp7_im_im_a2 0 x7_im_a2 1.6234265289688375e-10
Cx8_re_a2 x8_re_a2 0 1.0
Gx8_re_a2 0 x8_re_a2 p2 0 0.1414213562373095
Fx8_re_a2 0 x8_re_a2 V2 7.0710678118654755
Rp8_re_re_a2 0 x8_re_a2 1.4083143320865588e-10
Gp8_re_im_a2 0 x8_re_a2 x8_im_a2 0 175562128496.72046
Cx8_im_a2 x8_im_a2 0 1.0
Gp8_im_re_a2 0 x8_im_a2 x8_re_a2 0 -175562128496.72046
Rp8_im_im_a2 0 x8_im_a2 1.4083143320865588e-10
Cx9_re_a2 x9_re_a2 0 1.0
Gx9_re_a2 0 x9_re_a2 p2 0 0.1414213562373095
Fx9_re_a2 0 x9_re_a2 V2 7.0710678118654755
Rp9_re_re_a2 0 x9_re_a2 1.715215055825635e-10
Gp9_re_im_a2 0 x9_re_a2 x9_im_a2 0 170388268279.49786
Cx9_im_a2 x9_im_a2 0 1.0
Gp9_im_re_a2 0 x9_im_a2 x9_re_a2 0 -170388268279.49786
Rp9_im_im_a2 0 x9_im_a2 1.715215055825635e-10
Cx10_re_a2 x10_re_a2 0 1.0
Gx10_re_a2 0 x10_re_a2 p2 0 0.1414213562373095
Fx10_re_a2 0 x10_re_a2 V2 7.0710678118654755
Rp10_re_re_a2 0 x10_re_a2 1.279330633293622e-09
Gp10_re_im_a2 0 x10_re_a2 x10_im_a2 0 138925213075.38348
Cx10_im_a2 x10_im_a2 0 1.0
Gp10_im_re_a2 0 x10_im_a2 x10_re_a2 0 -138925213075.38348
Rp10_im_im_a2 0 x10_im_a2 1.279330633293622e-09
Cx11_re_a2 x11_re_a2 0 1.0
Gx11_re_a2 0 x11_re_a2 p2 0 0.1414213562373095
Fx11_re_a2 0 x11_re_a2 V2 7.0710678118654755
Rp11_re_re_a2 0 x11_re_a2 3.9059155840864643e-10
Gp11_re_im_a2 0 x11_re_a2 x11_im_a2 0 139719166370.31833
Cx11_im_a2 x11_im_a2 0 1.0
Gp11_im_re_a2 0 x11_im_a2 x11_re_a2 0 -139719166370.31833
Rp11_im_im_a2 0 x11_im_a2 3.9059155840864643e-10
Cx12_re_a2 x12_re_a2 0 1.0
Gx12_re_a2 0 x12_re_a2 p2 0 0.1414213562373095
Fx12_re_a2 0 x12_re_a2 V2 7.0710678118654755
Rp12_re_re_a2 0 x12_re_a2 1.049749481959773e-10
Gp12_re_im_a2 0 x12_re_a2 x12_im_a2 0 162806930635.2914
Cx12_im_a2 x12_im_a2 0 1.0
Gp12_im_re_a2 0 x12_im_a2 x12_re_a2 0 -162806930635.2914
Rp12_im_im_a2 0 x12_im_a2 1.049749481959773e-10
Cx13_re_a2 x13_re_a2 0 1.0
Gx13_re_a2 0 x13_re_a2 p2 0 0.1414213562373095
Fx13_re_a2 0 x13_re_a2 V2 7.0710678118654755
Rp13_re_re_a2 0 x13_re_a2 1.731638893406368e-10
Gp13_re_im_a2 0 x13_re_a2 x13_im_a2 0 161735038737.64923
Cx13_im_a2 x13_im_a2 0 1.0
Gp13_im_re_a2 0 x13_im_a2 x13_re_a2 0 -161735038737.64923
Rp13_im_im_a2 0 x13_im_a2 1.731638893406368e-10
Cx14_re_a2 x14_re_a2 0 1.0
Gx14_re_a2 0 x14_re_a2 p2 0 0.1414213562373095
Fx14_re_a2 0 x14_re_a2 V2 7.0710678118654755
Rp14_re_re_a2 0 x14_re_a2 1.5904302621228683e-10
Gp14_re_im_a2 0 x14_re_a2 x14_im_a2 0 154094455422.17636
Cx14_im_a2 x14_im_a2 0 1.0
Gp14_im_re_a2 0 x14_im_a2 x14_re_a2 0 -154094455422.17636
Rp14_im_im_a2 0 x14_im_a2 1.5904302621228683e-10
Cx15_re_a2 x15_re_a2 0 1.0
Gx15_re_a2 0 x15_re_a2 p2 0 0.1414213562373095
Fx15_re_a2 0 x15_re_a2 V2 7.0710678118654755
Rp15_re_re_a2 0 x15_re_a2 1.5963175233460748e-10
Gp15_re_im_a2 0 x15_re_a2 x15_im_a2 0 151958412904.65485
Cx15_im_a2 x15_im_a2 0 1.0
Gp15_im_re_a2 0 x15_im_a2 x15_re_a2 0 -151958412904.65485
Rp15_im_im_a2 0 x15_im_a2 1.5963175233460748e-10
Cx16_re_a2 x16_re_a2 0 1.0
Gx16_re_a2 0 x16_re_a2 p2 0 0.1414213562373095
Fx16_re_a2 0 x16_re_a2 V2 7.0710678118654755
Rp16_re_re_a2 0 x16_re_a2 4.085517959442536e-10
Gp16_re_im_a2 0 x16_re_a2 x16_im_a2 0 150304807574.39594
Cx16_im_a2 x16_im_a2 0 1.0
Gp16_im_re_a2 0 x16_im_a2 x16_re_a2 0 -150304807574.39594
Rp16_im_im_a2 0 x16_im_a2 4.085517959442536e-10
Cx17_re_a2 x17_re_a2 0 1.0
Gx17_re_a2 0 x17_re_a2 p2 0 0.1414213562373095
Fx17_re_a2 0 x17_re_a2 V2 7.0710678118654755
Rp17_re_re_a2 0 x17_re_a2 3.8552133160375805e-10
Gp17_re_im_a2 0 x17_re_a2 x17_im_a2 0 150713612315.05786
Cx17_im_a2 x17_im_a2 0 1.0
Gp17_im_re_a2 0 x17_im_a2 x17_re_a2 0 -150713612315.05786
Rp17_im_im_a2 0 x17_im_a2 3.8552133160375805e-10
.ENDS s_equivalent
