* EQUIVALENT CIRCUIT FOR VECTOR FITTED S-MATRIX
* Created using scikit-rf vectorFitting.py

.SUBCKT s_equivalent p1 p2 p3 p4 p5 p6 p7 p8 p9 p10 p11 p12 p13 p14 p15 p16 p17 p18

* Port network for port 1
R_ref_1 p1 a1 50.0
H_b_1 a1 0 V_c_1 14.142135623730951
* Differential incident wave a sources for transfer from port 1
H_p_1 nt_p_1 nts_p_1 H_b_1 3.5355339059327378
E_p_1 nts_p_1 0 p1 0 0.07071067811865475
E_n_1 0 nt_n_1 nt_p_1 0 1
* Current sensor on center node for transfer to port 1
V_c_1 nt_c_1 0 0
* Transfer network from port 1 to port 1
R1_1 nt_p_1 nt_c_1 0.0007564900050830436
X1 nt_p_1 nt_c_1 rl_admittance res=6.713812060922877e+16 ind=0.01239433452121846
X2 nt_n_1 nt_c_1 rl_admittance res=0.00045787217518182793 ind=2.0503953265122565e-14
X3 nt_p_1 nt_c_1 rl_admittance res=0.00054254751817662 ind=7.679384261163742e-14
X4 nt_p_1 nt_c_1 rl_admittance res=0.0005564228350387422 ind=3.0785512135842906e-13
X5 nt_n_1 nt_c_1 rl_admittance res=0.0005055304090704312 ind=1.4305226916553906e-13
X6 nt_n_1 nt_c_1 rl_admittance res=0.00047272890640632993 ind=8.643258284073119e-13
* Transfer network from port 2 to port 1
R1_2 nt_n_2 nt_c_1 0.003124999999999963
X7 nt_n_2 nt_c_1 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X8 nt_p_2 nt_c_1 rl_admittance res=187800143092.54297 ind=8.409869753766284
X9 nt_p_2 nt_c_1 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X10 nt_p_2 nt_c_1 rl_admittance res=63732557064.23586 ind=35.261662271871394
X11 nt_n_2 nt_c_1 rl_admittance res=112799484372.98152 ind=31.919389834390056
X12 nt_n_2 nt_c_1 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 3 to port 1
R1_3 nt_n_3 nt_c_1 0.003124999999999963
X13 nt_n_3 nt_c_1 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X14 nt_p_3 nt_c_1 rl_admittance res=187800143092.54297 ind=8.409869753766284
X15 nt_p_3 nt_c_1 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X16 nt_p_3 nt_c_1 rl_admittance res=63732557064.23586 ind=35.261662271871394
X17 nt_n_3 nt_c_1 rl_admittance res=112799484372.98152 ind=31.919389834390056
X18 nt_n_3 nt_c_1 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 4 to port 1
R1_4 nt_n_4 nt_c_1 0.003124999999999963
X19 nt_n_4 nt_c_1 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X20 nt_p_4 nt_c_1 rl_admittance res=187800143092.54297 ind=8.409869753766284
X21 nt_p_4 nt_c_1 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X22 nt_p_4 nt_c_1 rl_admittance res=63732557064.23586 ind=35.261662271871394
X23 nt_n_4 nt_c_1 rl_admittance res=112799484372.98152 ind=31.919389834390056
X24 nt_n_4 nt_c_1 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 5 to port 1
R1_5 nt_n_5 nt_c_1 0.003124999999999963
X25 nt_n_5 nt_c_1 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X26 nt_p_5 nt_c_1 rl_admittance res=187800143092.54297 ind=8.409869753766284
X27 nt_p_5 nt_c_1 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X28 nt_p_5 nt_c_1 rl_admittance res=63732557064.23586 ind=35.261662271871394
X29 nt_n_5 nt_c_1 rl_admittance res=112799484372.98152 ind=31.919389834390056
X30 nt_n_5 nt_c_1 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 6 to port 1
R1_6 nt_n_6 nt_c_1 0.003124999999999963
X31 nt_n_6 nt_c_1 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X32 nt_p_6 nt_c_1 rl_admittance res=187800143092.54297 ind=8.409869753766284
X33 nt_p_6 nt_c_1 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X34 nt_p_6 nt_c_1 rl_admittance res=63732557064.23586 ind=35.261662271871394
X35 nt_n_6 nt_c_1 rl_admittance res=112799484372.98152 ind=31.919389834390056
X36 nt_n_6 nt_c_1 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 7 to port 1
R1_7 nt_n_7 nt_c_1 0.003124999999999963
X37 nt_n_7 nt_c_1 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X38 nt_p_7 nt_c_1 rl_admittance res=187800143092.54297 ind=8.409869753766284
X39 nt_p_7 nt_c_1 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X40 nt_p_7 nt_c_1 rl_admittance res=63732557064.23586 ind=35.261662271871394
X41 nt_n_7 nt_c_1 rl_admittance res=112799484372.98152 ind=31.919389834390056
X42 nt_n_7 nt_c_1 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 8 to port 1
R1_8 nt_n_8 nt_c_1 0.003124999999999963
X43 nt_n_8 nt_c_1 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X44 nt_p_8 nt_c_1 rl_admittance res=187800143092.54297 ind=8.409869753766284
X45 nt_p_8 nt_c_1 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X46 nt_p_8 nt_c_1 rl_admittance res=63732557064.23586 ind=35.261662271871394
X47 nt_n_8 nt_c_1 rl_admittance res=112799484372.98152 ind=31.919389834390056
X48 nt_n_8 nt_c_1 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 9 to port 1
R1_9 nt_n_9 nt_c_1 0.003124999999999963
X49 nt_n_9 nt_c_1 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X50 nt_p_9 nt_c_1 rl_admittance res=187800143092.54297 ind=8.409869753766284
X51 nt_p_9 nt_c_1 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X52 nt_p_9 nt_c_1 rl_admittance res=63732557064.23586 ind=35.261662271871394
X53 nt_n_9 nt_c_1 rl_admittance res=112799484372.98152 ind=31.919389834390056
X54 nt_n_9 nt_c_1 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 10 to port 1
R1_10 nt_n_10 nt_c_1 0.003124999999999963
X55 nt_n_10 nt_c_1 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X56 nt_p_10 nt_c_1 rl_admittance res=187800143092.54297 ind=8.409869753766284
X57 nt_p_10 nt_c_1 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X58 nt_p_10 nt_c_1 rl_admittance res=63732557064.23586 ind=35.261662271871394
X59 nt_n_10 nt_c_1 rl_admittance res=112799484372.98152 ind=31.919389834390056
X60 nt_n_10 nt_c_1 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 11 to port 1
R1_11 nt_n_11 nt_c_1 0.003124999999999963
X61 nt_n_11 nt_c_1 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X62 nt_p_11 nt_c_1 rl_admittance res=187800143092.54297 ind=8.409869753766284
X63 nt_p_11 nt_c_1 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X64 nt_p_11 nt_c_1 rl_admittance res=63732557064.23586 ind=35.261662271871394
X65 nt_n_11 nt_c_1 rl_admittance res=112799484372.98152 ind=31.919389834390056
X66 nt_n_11 nt_c_1 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 12 to port 1
R1_12 nt_n_12 nt_c_1 0.003124999999999963
X67 nt_n_12 nt_c_1 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X68 nt_p_12 nt_c_1 rl_admittance res=187800143092.54297 ind=8.409869753766284
X69 nt_p_12 nt_c_1 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X70 nt_p_12 nt_c_1 rl_admittance res=63732557064.23586 ind=35.261662271871394
X71 nt_n_12 nt_c_1 rl_admittance res=112799484372.98152 ind=31.919389834390056
X72 nt_n_12 nt_c_1 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 13 to port 1
R1_13 nt_n_13 nt_c_1 0.003124999999999963
X73 nt_n_13 nt_c_1 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X74 nt_p_13 nt_c_1 rl_admittance res=187800143092.54297 ind=8.409869753766284
X75 nt_p_13 nt_c_1 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X76 nt_p_13 nt_c_1 rl_admittance res=63732557064.23586 ind=35.261662271871394
X77 nt_n_13 nt_c_1 rl_admittance res=112799484372.98152 ind=31.919389834390056
X78 nt_n_13 nt_c_1 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 14 to port 1
R1_14 nt_n_14 nt_c_1 0.003124999999999963
X79 nt_n_14 nt_c_1 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X80 nt_p_14 nt_c_1 rl_admittance res=187800143092.54297 ind=8.409869753766284
X81 nt_p_14 nt_c_1 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X82 nt_p_14 nt_c_1 rl_admittance res=63732557064.23586 ind=35.261662271871394
X83 nt_n_14 nt_c_1 rl_admittance res=112799484372.98152 ind=31.919389834390056
X84 nt_n_14 nt_c_1 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 15 to port 1
R1_15 nt_n_15 nt_c_1 0.003124999999999963
X85 nt_n_15 nt_c_1 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X86 nt_p_15 nt_c_1 rl_admittance res=187800143092.54297 ind=8.409869753766284
X87 nt_p_15 nt_c_1 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X88 nt_p_15 nt_c_1 rl_admittance res=63732557064.23586 ind=35.261662271871394
X89 nt_n_15 nt_c_1 rl_admittance res=112799484372.98152 ind=31.919389834390056
X90 nt_n_15 nt_c_1 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 16 to port 1
R1_16 nt_n_16 nt_c_1 0.003124999999999963
X91 nt_n_16 nt_c_1 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X92 nt_p_16 nt_c_1 rl_admittance res=187800143092.54297 ind=8.409869753766284
X93 nt_p_16 nt_c_1 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X94 nt_p_16 nt_c_1 rl_admittance res=63732557064.23586 ind=35.261662271871394
X95 nt_n_16 nt_c_1 rl_admittance res=112799484372.98152 ind=31.919389834390056
X96 nt_n_16 nt_c_1 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 17 to port 1
R1_17 nt_n_17 nt_c_1 0.003124999999999963
X97 nt_n_17 nt_c_1 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X98 nt_p_17 nt_c_1 rl_admittance res=187800143092.54297 ind=8.409869753766284
X99 nt_p_17 nt_c_1 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X100 nt_p_17 nt_c_1 rl_admittance res=63732557064.23586 ind=35.261662271871394
X101 nt_n_17 nt_c_1 rl_admittance res=112799484372.98152 ind=31.919389834390056
X102 nt_n_17 nt_c_1 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 18 to port 1
R1_18 nt_n_18 nt_c_1 0.003124999999999963
X103 nt_n_18 nt_c_1 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X104 nt_p_18 nt_c_1 rl_admittance res=187800143092.54297 ind=8.409869753766284
X105 nt_p_18 nt_c_1 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X106 nt_p_18 nt_c_1 rl_admittance res=63732557064.23586 ind=35.261662271871394
X107 nt_n_18 nt_c_1 rl_admittance res=112799484372.98152 ind=31.919389834390056
X108 nt_n_18 nt_c_1 rl_admittance res=51262611157.92125 ind=93.72728905498322

* Port network for port 2
R_ref_2 p2 a2 50.0
H_b_2 a2 0 V_c_2 14.142135623730951
* Differential incident wave a sources for transfer from port 2
H_p_2 nt_p_2 nts_p_2 H_b_2 3.5355339059327378
E_p_2 nts_p_2 0 p2 0 0.07071067811865475
E_n_2 0 nt_n_2 nt_p_2 0 1
* Current sensor on center node for transfer to port 2
V_c_2 nt_c_2 0 0
* Transfer network from port 1 to port 2
R2_1 nt_n_1 nt_c_2 0.003124999999999963
X109 nt_n_1 nt_c_2 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X110 nt_p_1 nt_c_2 rl_admittance res=187800143092.54297 ind=8.409869753766284
X111 nt_p_1 nt_c_2 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X112 nt_p_1 nt_c_2 rl_admittance res=63732557064.23586 ind=35.261662271871394
X113 nt_n_1 nt_c_2 rl_admittance res=112799484372.98152 ind=31.919389834390056
X114 nt_n_1 nt_c_2 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 2 to port 2
R2_2 nt_p_2 nt_c_2 0.0007564900050830436
X115 nt_p_2 nt_c_2 rl_admittance res=6.713812060922877e+16 ind=0.01239433452121846
X116 nt_n_2 nt_c_2 rl_admittance res=0.00045787217518182793 ind=2.0503953265122565e-14
X117 nt_p_2 nt_c_2 rl_admittance res=0.00054254751817662 ind=7.679384261163742e-14
X118 nt_p_2 nt_c_2 rl_admittance res=0.0005564228350387422 ind=3.0785512135842906e-13
X119 nt_n_2 nt_c_2 rl_admittance res=0.0005055304090704312 ind=1.4305226916553906e-13
X120 nt_n_2 nt_c_2 rl_admittance res=0.00047272890640632993 ind=8.643258284073119e-13
* Transfer network from port 3 to port 2
R2_3 nt_n_3 nt_c_2 0.003124999999999963
X121 nt_n_3 nt_c_2 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X122 nt_p_3 nt_c_2 rl_admittance res=187800143092.54297 ind=8.409869753766284
X123 nt_p_3 nt_c_2 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X124 nt_p_3 nt_c_2 rl_admittance res=63732557064.23586 ind=35.261662271871394
X125 nt_n_3 nt_c_2 rl_admittance res=112799484372.98152 ind=31.919389834390056
X126 nt_n_3 nt_c_2 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 4 to port 2
R2_4 nt_n_4 nt_c_2 0.003124999999999963
X127 nt_n_4 nt_c_2 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X128 nt_p_4 nt_c_2 rl_admittance res=187800143092.54297 ind=8.409869753766284
X129 nt_p_4 nt_c_2 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X130 nt_p_4 nt_c_2 rl_admittance res=63732557064.23586 ind=35.261662271871394
X131 nt_n_4 nt_c_2 rl_admittance res=112799484372.98152 ind=31.919389834390056
X132 nt_n_4 nt_c_2 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 5 to port 2
R2_5 nt_n_5 nt_c_2 0.003124999999999963
X133 nt_n_5 nt_c_2 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X134 nt_p_5 nt_c_2 rl_admittance res=187800143092.54297 ind=8.409869753766284
X135 nt_p_5 nt_c_2 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X136 nt_p_5 nt_c_2 rl_admittance res=63732557064.23586 ind=35.261662271871394
X137 nt_n_5 nt_c_2 rl_admittance res=112799484372.98152 ind=31.919389834390056
X138 nt_n_5 nt_c_2 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 6 to port 2
R2_6 nt_n_6 nt_c_2 0.003124999999999963
X139 nt_n_6 nt_c_2 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X140 nt_p_6 nt_c_2 rl_admittance res=187800143092.54297 ind=8.409869753766284
X141 nt_p_6 nt_c_2 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X142 nt_p_6 nt_c_2 rl_admittance res=63732557064.23586 ind=35.261662271871394
X143 nt_n_6 nt_c_2 rl_admittance res=112799484372.98152 ind=31.919389834390056
X144 nt_n_6 nt_c_2 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 7 to port 2
R2_7 nt_n_7 nt_c_2 0.003124999999999963
X145 nt_n_7 nt_c_2 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X146 nt_p_7 nt_c_2 rl_admittance res=187800143092.54297 ind=8.409869753766284
X147 nt_p_7 nt_c_2 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X148 nt_p_7 nt_c_2 rl_admittance res=63732557064.23586 ind=35.261662271871394
X149 nt_n_7 nt_c_2 rl_admittance res=112799484372.98152 ind=31.919389834390056
X150 nt_n_7 nt_c_2 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 8 to port 2
R2_8 nt_n_8 nt_c_2 0.003124999999999963
X151 nt_n_8 nt_c_2 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X152 nt_p_8 nt_c_2 rl_admittance res=187800143092.54297 ind=8.409869753766284
X153 nt_p_8 nt_c_2 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X154 nt_p_8 nt_c_2 rl_admittance res=63732557064.23586 ind=35.261662271871394
X155 nt_n_8 nt_c_2 rl_admittance res=112799484372.98152 ind=31.919389834390056
X156 nt_n_8 nt_c_2 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 9 to port 2
R2_9 nt_n_9 nt_c_2 0.003124999999999963
X157 nt_n_9 nt_c_2 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X158 nt_p_9 nt_c_2 rl_admittance res=187800143092.54297 ind=8.409869753766284
X159 nt_p_9 nt_c_2 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X160 nt_p_9 nt_c_2 rl_admittance res=63732557064.23586 ind=35.261662271871394
X161 nt_n_9 nt_c_2 rl_admittance res=112799484372.98152 ind=31.919389834390056
X162 nt_n_9 nt_c_2 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 10 to port 2
R2_10 nt_n_10 nt_c_2 0.003124999999999963
X163 nt_n_10 nt_c_2 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X164 nt_p_10 nt_c_2 rl_admittance res=187800143092.54297 ind=8.409869753766284
X165 nt_p_10 nt_c_2 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X166 nt_p_10 nt_c_2 rl_admittance res=63732557064.23586 ind=35.261662271871394
X167 nt_n_10 nt_c_2 rl_admittance res=112799484372.98152 ind=31.919389834390056
X168 nt_n_10 nt_c_2 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 11 to port 2
R2_11 nt_n_11 nt_c_2 0.003124999999999963
X169 nt_n_11 nt_c_2 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X170 nt_p_11 nt_c_2 rl_admittance res=187800143092.54297 ind=8.409869753766284
X171 nt_p_11 nt_c_2 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X172 nt_p_11 nt_c_2 rl_admittance res=63732557064.23586 ind=35.261662271871394
X173 nt_n_11 nt_c_2 rl_admittance res=112799484372.98152 ind=31.919389834390056
X174 nt_n_11 nt_c_2 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 12 to port 2
R2_12 nt_n_12 nt_c_2 0.003124999999999963
X175 nt_n_12 nt_c_2 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X176 nt_p_12 nt_c_2 rl_admittance res=187800143092.54297 ind=8.409869753766284
X177 nt_p_12 nt_c_2 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X178 nt_p_12 nt_c_2 rl_admittance res=63732557064.23586 ind=35.261662271871394
X179 nt_n_12 nt_c_2 rl_admittance res=112799484372.98152 ind=31.919389834390056
X180 nt_n_12 nt_c_2 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 13 to port 2
R2_13 nt_n_13 nt_c_2 0.003124999999999963
X181 nt_n_13 nt_c_2 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X182 nt_p_13 nt_c_2 rl_admittance res=187800143092.54297 ind=8.409869753766284
X183 nt_p_13 nt_c_2 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X184 nt_p_13 nt_c_2 rl_admittance res=63732557064.23586 ind=35.261662271871394
X185 nt_n_13 nt_c_2 rl_admittance res=112799484372.98152 ind=31.919389834390056
X186 nt_n_13 nt_c_2 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 14 to port 2
R2_14 nt_n_14 nt_c_2 0.003124999999999963
X187 nt_n_14 nt_c_2 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X188 nt_p_14 nt_c_2 rl_admittance res=187800143092.54297 ind=8.409869753766284
X189 nt_p_14 nt_c_2 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X190 nt_p_14 nt_c_2 rl_admittance res=63732557064.23586 ind=35.261662271871394
X191 nt_n_14 nt_c_2 rl_admittance res=112799484372.98152 ind=31.919389834390056
X192 nt_n_14 nt_c_2 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 15 to port 2
R2_15 nt_n_15 nt_c_2 0.003124999999999963
X193 nt_n_15 nt_c_2 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X194 nt_p_15 nt_c_2 rl_admittance res=187800143092.54297 ind=8.409869753766284
X195 nt_p_15 nt_c_2 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X196 nt_p_15 nt_c_2 rl_admittance res=63732557064.23586 ind=35.261662271871394
X197 nt_n_15 nt_c_2 rl_admittance res=112799484372.98152 ind=31.919389834390056
X198 nt_n_15 nt_c_2 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 16 to port 2
R2_16 nt_n_16 nt_c_2 0.003124999999999963
X199 nt_n_16 nt_c_2 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X200 nt_p_16 nt_c_2 rl_admittance res=187800143092.54297 ind=8.409869753766284
X201 nt_p_16 nt_c_2 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X202 nt_p_16 nt_c_2 rl_admittance res=63732557064.23586 ind=35.261662271871394
X203 nt_n_16 nt_c_2 rl_admittance res=112799484372.98152 ind=31.919389834390056
X204 nt_n_16 nt_c_2 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 17 to port 2
R2_17 nt_n_17 nt_c_2 0.003124999999999963
X205 nt_n_17 nt_c_2 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X206 nt_p_17 nt_c_2 rl_admittance res=187800143092.54297 ind=8.409869753766284
X207 nt_p_17 nt_c_2 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X208 nt_p_17 nt_c_2 rl_admittance res=63732557064.23586 ind=35.261662271871394
X209 nt_n_17 nt_c_2 rl_admittance res=112799484372.98152 ind=31.919389834390056
X210 nt_n_17 nt_c_2 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 18 to port 2
R2_18 nt_n_18 nt_c_2 0.003124999999999963
X211 nt_n_18 nt_c_2 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X212 nt_p_18 nt_c_2 rl_admittance res=187800143092.54297 ind=8.409869753766284
X213 nt_p_18 nt_c_2 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X214 nt_p_18 nt_c_2 rl_admittance res=63732557064.23586 ind=35.261662271871394
X215 nt_n_18 nt_c_2 rl_admittance res=112799484372.98152 ind=31.919389834390056
X216 nt_n_18 nt_c_2 rl_admittance res=51262611157.92125 ind=93.72728905498322

* Port network for port 3
R_ref_3 p3 a3 50.0
H_b_3 a3 0 V_c_3 14.142135623730951
* Differential incident wave a sources for transfer from port 3
H_p_3 nt_p_3 nts_p_3 H_b_3 3.5355339059327378
E_p_3 nts_p_3 0 p3 0 0.07071067811865475
E_n_3 0 nt_n_3 nt_p_3 0 1
* Current sensor on center node for transfer to port 3
V_c_3 nt_c_3 0 0
* Transfer network from port 1 to port 3
R3_1 nt_n_1 nt_c_3 0.003124999999999963
X217 nt_n_1 nt_c_3 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X218 nt_p_1 nt_c_3 rl_admittance res=187800143092.54297 ind=8.409869753766284
X219 nt_p_1 nt_c_3 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X220 nt_p_1 nt_c_3 rl_admittance res=63732557064.23586 ind=35.261662271871394
X221 nt_n_1 nt_c_3 rl_admittance res=112799484372.98152 ind=31.919389834390056
X222 nt_n_1 nt_c_3 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 2 to port 3
R3_2 nt_n_2 nt_c_3 0.003124999999999963
X223 nt_n_2 nt_c_3 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X224 nt_p_2 nt_c_3 rl_admittance res=187800143092.54297 ind=8.409869753766284
X225 nt_p_2 nt_c_3 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X226 nt_p_2 nt_c_3 rl_admittance res=63732557064.23586 ind=35.261662271871394
X227 nt_n_2 nt_c_3 rl_admittance res=112799484372.98152 ind=31.919389834390056
X228 nt_n_2 nt_c_3 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 3 to port 3
R3_3 nt_p_3 nt_c_3 0.0007564900050830436
X229 nt_p_3 nt_c_3 rl_admittance res=6.713812060922877e+16 ind=0.01239433452121846
X230 nt_n_3 nt_c_3 rl_admittance res=0.00045787217518182793 ind=2.0503953265122565e-14
X231 nt_p_3 nt_c_3 rl_admittance res=0.00054254751817662 ind=7.679384261163742e-14
X232 nt_p_3 nt_c_3 rl_admittance res=0.0005564228350387422 ind=3.0785512135842906e-13
X233 nt_n_3 nt_c_3 rl_admittance res=0.0005055304090704312 ind=1.4305226916553906e-13
X234 nt_n_3 nt_c_3 rl_admittance res=0.00047272890640632993 ind=8.643258284073119e-13
* Transfer network from port 4 to port 3
R3_4 nt_n_4 nt_c_3 0.003124999999999963
X235 nt_n_4 nt_c_3 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X236 nt_p_4 nt_c_3 rl_admittance res=187800143092.54297 ind=8.409869753766284
X237 nt_p_4 nt_c_3 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X238 nt_p_4 nt_c_3 rl_admittance res=63732557064.23586 ind=35.261662271871394
X239 nt_n_4 nt_c_3 rl_admittance res=112799484372.98152 ind=31.919389834390056
X240 nt_n_4 nt_c_3 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 5 to port 3
R3_5 nt_n_5 nt_c_3 0.003124999999999963
X241 nt_n_5 nt_c_3 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X242 nt_p_5 nt_c_3 rl_admittance res=187800143092.54297 ind=8.409869753766284
X243 nt_p_5 nt_c_3 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X244 nt_p_5 nt_c_3 rl_admittance res=63732557064.23586 ind=35.261662271871394
X245 nt_n_5 nt_c_3 rl_admittance res=112799484372.98152 ind=31.919389834390056
X246 nt_n_5 nt_c_3 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 6 to port 3
R3_6 nt_n_6 nt_c_3 0.003124999999999963
X247 nt_n_6 nt_c_3 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X248 nt_p_6 nt_c_3 rl_admittance res=187800143092.54297 ind=8.409869753766284
X249 nt_p_6 nt_c_3 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X250 nt_p_6 nt_c_3 rl_admittance res=63732557064.23586 ind=35.261662271871394
X251 nt_n_6 nt_c_3 rl_admittance res=112799484372.98152 ind=31.919389834390056
X252 nt_n_6 nt_c_3 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 7 to port 3
R3_7 nt_n_7 nt_c_3 0.003124999999999963
X253 nt_n_7 nt_c_3 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X254 nt_p_7 nt_c_3 rl_admittance res=187800143092.54297 ind=8.409869753766284
X255 nt_p_7 nt_c_3 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X256 nt_p_7 nt_c_3 rl_admittance res=63732557064.23586 ind=35.261662271871394
X257 nt_n_7 nt_c_3 rl_admittance res=112799484372.98152 ind=31.919389834390056
X258 nt_n_7 nt_c_3 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 8 to port 3
R3_8 nt_n_8 nt_c_3 0.003124999999999963
X259 nt_n_8 nt_c_3 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X260 nt_p_8 nt_c_3 rl_admittance res=187800143092.54297 ind=8.409869753766284
X261 nt_p_8 nt_c_3 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X262 nt_p_8 nt_c_3 rl_admittance res=63732557064.23586 ind=35.261662271871394
X263 nt_n_8 nt_c_3 rl_admittance res=112799484372.98152 ind=31.919389834390056
X264 nt_n_8 nt_c_3 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 9 to port 3
R3_9 nt_n_9 nt_c_3 0.003124999999999963
X265 nt_n_9 nt_c_3 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X266 nt_p_9 nt_c_3 rl_admittance res=187800143092.54297 ind=8.409869753766284
X267 nt_p_9 nt_c_3 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X268 nt_p_9 nt_c_3 rl_admittance res=63732557064.23586 ind=35.261662271871394
X269 nt_n_9 nt_c_3 rl_admittance res=112799484372.98152 ind=31.919389834390056
X270 nt_n_9 nt_c_3 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 10 to port 3
R3_10 nt_n_10 nt_c_3 0.003124999999999963
X271 nt_n_10 nt_c_3 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X272 nt_p_10 nt_c_3 rl_admittance res=187800143092.54297 ind=8.409869753766284
X273 nt_p_10 nt_c_3 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X274 nt_p_10 nt_c_3 rl_admittance res=63732557064.23586 ind=35.261662271871394
X275 nt_n_10 nt_c_3 rl_admittance res=112799484372.98152 ind=31.919389834390056
X276 nt_n_10 nt_c_3 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 11 to port 3
R3_11 nt_n_11 nt_c_3 0.003124999999999963
X277 nt_n_11 nt_c_3 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X278 nt_p_11 nt_c_3 rl_admittance res=187800143092.54297 ind=8.409869753766284
X279 nt_p_11 nt_c_3 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X280 nt_p_11 nt_c_3 rl_admittance res=63732557064.23586 ind=35.261662271871394
X281 nt_n_11 nt_c_3 rl_admittance res=112799484372.98152 ind=31.919389834390056
X282 nt_n_11 nt_c_3 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 12 to port 3
R3_12 nt_n_12 nt_c_3 0.003124999999999963
X283 nt_n_12 nt_c_3 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X284 nt_p_12 nt_c_3 rl_admittance res=187800143092.54297 ind=8.409869753766284
X285 nt_p_12 nt_c_3 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X286 nt_p_12 nt_c_3 rl_admittance res=63732557064.23586 ind=35.261662271871394
X287 nt_n_12 nt_c_3 rl_admittance res=112799484372.98152 ind=31.919389834390056
X288 nt_n_12 nt_c_3 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 13 to port 3
R3_13 nt_n_13 nt_c_3 0.003124999999999963
X289 nt_n_13 nt_c_3 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X290 nt_p_13 nt_c_3 rl_admittance res=187800143092.54297 ind=8.409869753766284
X291 nt_p_13 nt_c_3 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X292 nt_p_13 nt_c_3 rl_admittance res=63732557064.23586 ind=35.261662271871394
X293 nt_n_13 nt_c_3 rl_admittance res=112799484372.98152 ind=31.919389834390056
X294 nt_n_13 nt_c_3 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 14 to port 3
R3_14 nt_n_14 nt_c_3 0.003124999999999963
X295 nt_n_14 nt_c_3 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X296 nt_p_14 nt_c_3 rl_admittance res=187800143092.54297 ind=8.409869753766284
X297 nt_p_14 nt_c_3 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X298 nt_p_14 nt_c_3 rl_admittance res=63732557064.23586 ind=35.261662271871394
X299 nt_n_14 nt_c_3 rl_admittance res=112799484372.98152 ind=31.919389834390056
X300 nt_n_14 nt_c_3 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 15 to port 3
R3_15 nt_n_15 nt_c_3 0.003124999999999963
X301 nt_n_15 nt_c_3 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X302 nt_p_15 nt_c_3 rl_admittance res=187800143092.54297 ind=8.409869753766284
X303 nt_p_15 nt_c_3 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X304 nt_p_15 nt_c_3 rl_admittance res=63732557064.23586 ind=35.261662271871394
X305 nt_n_15 nt_c_3 rl_admittance res=112799484372.98152 ind=31.919389834390056
X306 nt_n_15 nt_c_3 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 16 to port 3
R3_16 nt_n_16 nt_c_3 0.003124999999999963
X307 nt_n_16 nt_c_3 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X308 nt_p_16 nt_c_3 rl_admittance res=187800143092.54297 ind=8.409869753766284
X309 nt_p_16 nt_c_3 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X310 nt_p_16 nt_c_3 rl_admittance res=63732557064.23586 ind=35.261662271871394
X311 nt_n_16 nt_c_3 rl_admittance res=112799484372.98152 ind=31.919389834390056
X312 nt_n_16 nt_c_3 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 17 to port 3
R3_17 nt_n_17 nt_c_3 0.003124999999999963
X313 nt_n_17 nt_c_3 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X314 nt_p_17 nt_c_3 rl_admittance res=187800143092.54297 ind=8.409869753766284
X315 nt_p_17 nt_c_3 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X316 nt_p_17 nt_c_3 rl_admittance res=63732557064.23586 ind=35.261662271871394
X317 nt_n_17 nt_c_3 rl_admittance res=112799484372.98152 ind=31.919389834390056
X318 nt_n_17 nt_c_3 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 18 to port 3
R3_18 nt_n_18 nt_c_3 0.003124999999999963
X319 nt_n_18 nt_c_3 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X320 nt_p_18 nt_c_3 rl_admittance res=187800143092.54297 ind=8.409869753766284
X321 nt_p_18 nt_c_3 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X322 nt_p_18 nt_c_3 rl_admittance res=63732557064.23586 ind=35.261662271871394
X323 nt_n_18 nt_c_3 rl_admittance res=112799484372.98152 ind=31.919389834390056
X324 nt_n_18 nt_c_3 rl_admittance res=51262611157.92125 ind=93.72728905498322

* Port network for port 4
R_ref_4 p4 a4 50.0
H_b_4 a4 0 V_c_4 14.142135623730951
* Differential incident wave a sources for transfer from port 4
H_p_4 nt_p_4 nts_p_4 H_b_4 3.5355339059327378
E_p_4 nts_p_4 0 p4 0 0.07071067811865475
E_n_4 0 nt_n_4 nt_p_4 0 1
* Current sensor on center node for transfer to port 4
V_c_4 nt_c_4 0 0
* Transfer network from port 1 to port 4
R4_1 nt_n_1 nt_c_4 0.003124999999999963
X325 nt_n_1 nt_c_4 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X326 nt_p_1 nt_c_4 rl_admittance res=187800143092.54297 ind=8.409869753766284
X327 nt_p_1 nt_c_4 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X328 nt_p_1 nt_c_4 rl_admittance res=63732557064.23586 ind=35.261662271871394
X329 nt_n_1 nt_c_4 rl_admittance res=112799484372.98152 ind=31.919389834390056
X330 nt_n_1 nt_c_4 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 2 to port 4
R4_2 nt_n_2 nt_c_4 0.003124999999999963
X331 nt_n_2 nt_c_4 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X332 nt_p_2 nt_c_4 rl_admittance res=187800143092.54297 ind=8.409869753766284
X333 nt_p_2 nt_c_4 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X334 nt_p_2 nt_c_4 rl_admittance res=63732557064.23586 ind=35.261662271871394
X335 nt_n_2 nt_c_4 rl_admittance res=112799484372.98152 ind=31.919389834390056
X336 nt_n_2 nt_c_4 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 3 to port 4
R4_3 nt_n_3 nt_c_4 0.003124999999999963
X337 nt_n_3 nt_c_4 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X338 nt_p_3 nt_c_4 rl_admittance res=187800143092.54297 ind=8.409869753766284
X339 nt_p_3 nt_c_4 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X340 nt_p_3 nt_c_4 rl_admittance res=63732557064.23586 ind=35.261662271871394
X341 nt_n_3 nt_c_4 rl_admittance res=112799484372.98152 ind=31.919389834390056
X342 nt_n_3 nt_c_4 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 4 to port 4
R4_4 nt_p_4 nt_c_4 0.0007564900050830436
X343 nt_p_4 nt_c_4 rl_admittance res=6.713812060922877e+16 ind=0.01239433452121846
X344 nt_n_4 nt_c_4 rl_admittance res=0.00045787217518182793 ind=2.0503953265122565e-14
X345 nt_p_4 nt_c_4 rl_admittance res=0.00054254751817662 ind=7.679384261163742e-14
X346 nt_p_4 nt_c_4 rl_admittance res=0.0005564228350387422 ind=3.0785512135842906e-13
X347 nt_n_4 nt_c_4 rl_admittance res=0.0005055304090704312 ind=1.4305226916553906e-13
X348 nt_n_4 nt_c_4 rl_admittance res=0.00047272890640632993 ind=8.643258284073119e-13
* Transfer network from port 5 to port 4
R4_5 nt_n_5 nt_c_4 0.003124999999999963
X349 nt_n_5 nt_c_4 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X350 nt_p_5 nt_c_4 rl_admittance res=187800143092.54297 ind=8.409869753766284
X351 nt_p_5 nt_c_4 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X352 nt_p_5 nt_c_4 rl_admittance res=63732557064.23586 ind=35.261662271871394
X353 nt_n_5 nt_c_4 rl_admittance res=112799484372.98152 ind=31.919389834390056
X354 nt_n_5 nt_c_4 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 6 to port 4
R4_6 nt_n_6 nt_c_4 0.003124999999999963
X355 nt_n_6 nt_c_4 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X356 nt_p_6 nt_c_4 rl_admittance res=187800143092.54297 ind=8.409869753766284
X357 nt_p_6 nt_c_4 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X358 nt_p_6 nt_c_4 rl_admittance res=63732557064.23586 ind=35.261662271871394
X359 nt_n_6 nt_c_4 rl_admittance res=112799484372.98152 ind=31.919389834390056
X360 nt_n_6 nt_c_4 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 7 to port 4
R4_7 nt_n_7 nt_c_4 0.003124999999999963
X361 nt_n_7 nt_c_4 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X362 nt_p_7 nt_c_4 rl_admittance res=187800143092.54297 ind=8.409869753766284
X363 nt_p_7 nt_c_4 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X364 nt_p_7 nt_c_4 rl_admittance res=63732557064.23586 ind=35.261662271871394
X365 nt_n_7 nt_c_4 rl_admittance res=112799484372.98152 ind=31.919389834390056
X366 nt_n_7 nt_c_4 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 8 to port 4
R4_8 nt_n_8 nt_c_4 0.003124999999999963
X367 nt_n_8 nt_c_4 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X368 nt_p_8 nt_c_4 rl_admittance res=187800143092.54297 ind=8.409869753766284
X369 nt_p_8 nt_c_4 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X370 nt_p_8 nt_c_4 rl_admittance res=63732557064.23586 ind=35.261662271871394
X371 nt_n_8 nt_c_4 rl_admittance res=112799484372.98152 ind=31.919389834390056
X372 nt_n_8 nt_c_4 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 9 to port 4
R4_9 nt_n_9 nt_c_4 0.003124999999999963
X373 nt_n_9 nt_c_4 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X374 nt_p_9 nt_c_4 rl_admittance res=187800143092.54297 ind=8.409869753766284
X375 nt_p_9 nt_c_4 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X376 nt_p_9 nt_c_4 rl_admittance res=63732557064.23586 ind=35.261662271871394
X377 nt_n_9 nt_c_4 rl_admittance res=112799484372.98152 ind=31.919389834390056
X378 nt_n_9 nt_c_4 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 10 to port 4
R4_10 nt_n_10 nt_c_4 0.003124999999999963
X379 nt_n_10 nt_c_4 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X380 nt_p_10 nt_c_4 rl_admittance res=187800143092.54297 ind=8.409869753766284
X381 nt_p_10 nt_c_4 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X382 nt_p_10 nt_c_4 rl_admittance res=63732557064.23586 ind=35.261662271871394
X383 nt_n_10 nt_c_4 rl_admittance res=112799484372.98152 ind=31.919389834390056
X384 nt_n_10 nt_c_4 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 11 to port 4
R4_11 nt_n_11 nt_c_4 0.003124999999999963
X385 nt_n_11 nt_c_4 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X386 nt_p_11 nt_c_4 rl_admittance res=187800143092.54297 ind=8.409869753766284
X387 nt_p_11 nt_c_4 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X388 nt_p_11 nt_c_4 rl_admittance res=63732557064.23586 ind=35.261662271871394
X389 nt_n_11 nt_c_4 rl_admittance res=112799484372.98152 ind=31.919389834390056
X390 nt_n_11 nt_c_4 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 12 to port 4
R4_12 nt_n_12 nt_c_4 0.003124999999999963
X391 nt_n_12 nt_c_4 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X392 nt_p_12 nt_c_4 rl_admittance res=187800143092.54297 ind=8.409869753766284
X393 nt_p_12 nt_c_4 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X394 nt_p_12 nt_c_4 rl_admittance res=63732557064.23586 ind=35.261662271871394
X395 nt_n_12 nt_c_4 rl_admittance res=112799484372.98152 ind=31.919389834390056
X396 nt_n_12 nt_c_4 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 13 to port 4
R4_13 nt_n_13 nt_c_4 0.003124999999999963
X397 nt_n_13 nt_c_4 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X398 nt_p_13 nt_c_4 rl_admittance res=187800143092.54297 ind=8.409869753766284
X399 nt_p_13 nt_c_4 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X400 nt_p_13 nt_c_4 rl_admittance res=63732557064.23586 ind=35.261662271871394
X401 nt_n_13 nt_c_4 rl_admittance res=112799484372.98152 ind=31.919389834390056
X402 nt_n_13 nt_c_4 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 14 to port 4
R4_14 nt_n_14 nt_c_4 0.003124999999999963
X403 nt_n_14 nt_c_4 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X404 nt_p_14 nt_c_4 rl_admittance res=187800143092.54297 ind=8.409869753766284
X405 nt_p_14 nt_c_4 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X406 nt_p_14 nt_c_4 rl_admittance res=63732557064.23586 ind=35.261662271871394
X407 nt_n_14 nt_c_4 rl_admittance res=112799484372.98152 ind=31.919389834390056
X408 nt_n_14 nt_c_4 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 15 to port 4
R4_15 nt_n_15 nt_c_4 0.003124999999999963
X409 nt_n_15 nt_c_4 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X410 nt_p_15 nt_c_4 rl_admittance res=187800143092.54297 ind=8.409869753766284
X411 nt_p_15 nt_c_4 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X412 nt_p_15 nt_c_4 rl_admittance res=63732557064.23586 ind=35.261662271871394
X413 nt_n_15 nt_c_4 rl_admittance res=112799484372.98152 ind=31.919389834390056
X414 nt_n_15 nt_c_4 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 16 to port 4
R4_16 nt_n_16 nt_c_4 0.003124999999999963
X415 nt_n_16 nt_c_4 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X416 nt_p_16 nt_c_4 rl_admittance res=187800143092.54297 ind=8.409869753766284
X417 nt_p_16 nt_c_4 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X418 nt_p_16 nt_c_4 rl_admittance res=63732557064.23586 ind=35.261662271871394
X419 nt_n_16 nt_c_4 rl_admittance res=112799484372.98152 ind=31.919389834390056
X420 nt_n_16 nt_c_4 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 17 to port 4
R4_17 nt_n_17 nt_c_4 0.003124999999999963
X421 nt_n_17 nt_c_4 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X422 nt_p_17 nt_c_4 rl_admittance res=187800143092.54297 ind=8.409869753766284
X423 nt_p_17 nt_c_4 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X424 nt_p_17 nt_c_4 rl_admittance res=63732557064.23586 ind=35.261662271871394
X425 nt_n_17 nt_c_4 rl_admittance res=112799484372.98152 ind=31.919389834390056
X426 nt_n_17 nt_c_4 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 18 to port 4
R4_18 nt_n_18 nt_c_4 0.003124999999999963
X427 nt_n_18 nt_c_4 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X428 nt_p_18 nt_c_4 rl_admittance res=187800143092.54297 ind=8.409869753766284
X429 nt_p_18 nt_c_4 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X430 nt_p_18 nt_c_4 rl_admittance res=63732557064.23586 ind=35.261662271871394
X431 nt_n_18 nt_c_4 rl_admittance res=112799484372.98152 ind=31.919389834390056
X432 nt_n_18 nt_c_4 rl_admittance res=51262611157.92125 ind=93.72728905498322

* Port network for port 5
R_ref_5 p5 a5 50.0
H_b_5 a5 0 V_c_5 14.142135623730951
* Differential incident wave a sources for transfer from port 5
H_p_5 nt_p_5 nts_p_5 H_b_5 3.5355339059327378
E_p_5 nts_p_5 0 p5 0 0.07071067811865475
E_n_5 0 nt_n_5 nt_p_5 0 1
* Current sensor on center node for transfer to port 5
V_c_5 nt_c_5 0 0
* Transfer network from port 1 to port 5
R5_1 nt_n_1 nt_c_5 0.003124999999999963
X433 nt_n_1 nt_c_5 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X434 nt_p_1 nt_c_5 rl_admittance res=187800143092.54297 ind=8.409869753766284
X435 nt_p_1 nt_c_5 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X436 nt_p_1 nt_c_5 rl_admittance res=63732557064.23586 ind=35.261662271871394
X437 nt_n_1 nt_c_5 rl_admittance res=112799484372.98152 ind=31.919389834390056
X438 nt_n_1 nt_c_5 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 2 to port 5
R5_2 nt_n_2 nt_c_5 0.003124999999999963
X439 nt_n_2 nt_c_5 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X440 nt_p_2 nt_c_5 rl_admittance res=187800143092.54297 ind=8.409869753766284
X441 nt_p_2 nt_c_5 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X442 nt_p_2 nt_c_5 rl_admittance res=63732557064.23586 ind=35.261662271871394
X443 nt_n_2 nt_c_5 rl_admittance res=112799484372.98152 ind=31.919389834390056
X444 nt_n_2 nt_c_5 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 3 to port 5
R5_3 nt_n_3 nt_c_5 0.003124999999999963
X445 nt_n_3 nt_c_5 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X446 nt_p_3 nt_c_5 rl_admittance res=187800143092.54297 ind=8.409869753766284
X447 nt_p_3 nt_c_5 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X448 nt_p_3 nt_c_5 rl_admittance res=63732557064.23586 ind=35.261662271871394
X449 nt_n_3 nt_c_5 rl_admittance res=112799484372.98152 ind=31.919389834390056
X450 nt_n_3 nt_c_5 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 4 to port 5
R5_4 nt_n_4 nt_c_5 0.003124999999999963
X451 nt_n_4 nt_c_5 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X452 nt_p_4 nt_c_5 rl_admittance res=187800143092.54297 ind=8.409869753766284
X453 nt_p_4 nt_c_5 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X454 nt_p_4 nt_c_5 rl_admittance res=63732557064.23586 ind=35.261662271871394
X455 nt_n_4 nt_c_5 rl_admittance res=112799484372.98152 ind=31.919389834390056
X456 nt_n_4 nt_c_5 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 5 to port 5
R5_5 nt_p_5 nt_c_5 0.0007564900050830436
X457 nt_p_5 nt_c_5 rl_admittance res=6.713812060922877e+16 ind=0.01239433452121846
X458 nt_n_5 nt_c_5 rl_admittance res=0.00045787217518182793 ind=2.0503953265122565e-14
X459 nt_p_5 nt_c_5 rl_admittance res=0.00054254751817662 ind=7.679384261163742e-14
X460 nt_p_5 nt_c_5 rl_admittance res=0.0005564228350387422 ind=3.0785512135842906e-13
X461 nt_n_5 nt_c_5 rl_admittance res=0.0005055304090704312 ind=1.4305226916553906e-13
X462 nt_n_5 nt_c_5 rl_admittance res=0.00047272890640632993 ind=8.643258284073119e-13
* Transfer network from port 6 to port 5
R5_6 nt_n_6 nt_c_5 0.003124999999999963
X463 nt_n_6 nt_c_5 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X464 nt_p_6 nt_c_5 rl_admittance res=187800143092.54297 ind=8.409869753766284
X465 nt_p_6 nt_c_5 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X466 nt_p_6 nt_c_5 rl_admittance res=63732557064.23586 ind=35.261662271871394
X467 nt_n_6 nt_c_5 rl_admittance res=112799484372.98152 ind=31.919389834390056
X468 nt_n_6 nt_c_5 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 7 to port 5
R5_7 nt_n_7 nt_c_5 0.003124999999999963
X469 nt_n_7 nt_c_5 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X470 nt_p_7 nt_c_5 rl_admittance res=187800143092.54297 ind=8.409869753766284
X471 nt_p_7 nt_c_5 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X472 nt_p_7 nt_c_5 rl_admittance res=63732557064.23586 ind=35.261662271871394
X473 nt_n_7 nt_c_5 rl_admittance res=112799484372.98152 ind=31.919389834390056
X474 nt_n_7 nt_c_5 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 8 to port 5
R5_8 nt_n_8 nt_c_5 0.003124999999999963
X475 nt_n_8 nt_c_5 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X476 nt_p_8 nt_c_5 rl_admittance res=187800143092.54297 ind=8.409869753766284
X477 nt_p_8 nt_c_5 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X478 nt_p_8 nt_c_5 rl_admittance res=63732557064.23586 ind=35.261662271871394
X479 nt_n_8 nt_c_5 rl_admittance res=112799484372.98152 ind=31.919389834390056
X480 nt_n_8 nt_c_5 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 9 to port 5
R5_9 nt_n_9 nt_c_5 0.003124999999999963
X481 nt_n_9 nt_c_5 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X482 nt_p_9 nt_c_5 rl_admittance res=187800143092.54297 ind=8.409869753766284
X483 nt_p_9 nt_c_5 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X484 nt_p_9 nt_c_5 rl_admittance res=63732557064.23586 ind=35.261662271871394
X485 nt_n_9 nt_c_5 rl_admittance res=112799484372.98152 ind=31.919389834390056
X486 nt_n_9 nt_c_5 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 10 to port 5
R5_10 nt_n_10 nt_c_5 0.003124999999999963
X487 nt_n_10 nt_c_5 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X488 nt_p_10 nt_c_5 rl_admittance res=187800143092.54297 ind=8.409869753766284
X489 nt_p_10 nt_c_5 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X490 nt_p_10 nt_c_5 rl_admittance res=63732557064.23586 ind=35.261662271871394
X491 nt_n_10 nt_c_5 rl_admittance res=112799484372.98152 ind=31.919389834390056
X492 nt_n_10 nt_c_5 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 11 to port 5
R5_11 nt_n_11 nt_c_5 0.003124999999999963
X493 nt_n_11 nt_c_5 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X494 nt_p_11 nt_c_5 rl_admittance res=187800143092.54297 ind=8.409869753766284
X495 nt_p_11 nt_c_5 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X496 nt_p_11 nt_c_5 rl_admittance res=63732557064.23586 ind=35.261662271871394
X497 nt_n_11 nt_c_5 rl_admittance res=112799484372.98152 ind=31.919389834390056
X498 nt_n_11 nt_c_5 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 12 to port 5
R5_12 nt_n_12 nt_c_5 0.003124999999999963
X499 nt_n_12 nt_c_5 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X500 nt_p_12 nt_c_5 rl_admittance res=187800143092.54297 ind=8.409869753766284
X501 nt_p_12 nt_c_5 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X502 nt_p_12 nt_c_5 rl_admittance res=63732557064.23586 ind=35.261662271871394
X503 nt_n_12 nt_c_5 rl_admittance res=112799484372.98152 ind=31.919389834390056
X504 nt_n_12 nt_c_5 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 13 to port 5
R5_13 nt_n_13 nt_c_5 0.003124999999999963
X505 nt_n_13 nt_c_5 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X506 nt_p_13 nt_c_5 rl_admittance res=187800143092.54297 ind=8.409869753766284
X507 nt_p_13 nt_c_5 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X508 nt_p_13 nt_c_5 rl_admittance res=63732557064.23586 ind=35.261662271871394
X509 nt_n_13 nt_c_5 rl_admittance res=112799484372.98152 ind=31.919389834390056
X510 nt_n_13 nt_c_5 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 14 to port 5
R5_14 nt_n_14 nt_c_5 0.003124999999999963
X511 nt_n_14 nt_c_5 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X512 nt_p_14 nt_c_5 rl_admittance res=187800143092.54297 ind=8.409869753766284
X513 nt_p_14 nt_c_5 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X514 nt_p_14 nt_c_5 rl_admittance res=63732557064.23586 ind=35.261662271871394
X515 nt_n_14 nt_c_5 rl_admittance res=112799484372.98152 ind=31.919389834390056
X516 nt_n_14 nt_c_5 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 15 to port 5
R5_15 nt_n_15 nt_c_5 0.003124999999999963
X517 nt_n_15 nt_c_5 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X518 nt_p_15 nt_c_5 rl_admittance res=187800143092.54297 ind=8.409869753766284
X519 nt_p_15 nt_c_5 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X520 nt_p_15 nt_c_5 rl_admittance res=63732557064.23586 ind=35.261662271871394
X521 nt_n_15 nt_c_5 rl_admittance res=112799484372.98152 ind=31.919389834390056
X522 nt_n_15 nt_c_5 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 16 to port 5
R5_16 nt_n_16 nt_c_5 0.003124999999999963
X523 nt_n_16 nt_c_5 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X524 nt_p_16 nt_c_5 rl_admittance res=187800143092.54297 ind=8.409869753766284
X525 nt_p_16 nt_c_5 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X526 nt_p_16 nt_c_5 rl_admittance res=63732557064.23586 ind=35.261662271871394
X527 nt_n_16 nt_c_5 rl_admittance res=112799484372.98152 ind=31.919389834390056
X528 nt_n_16 nt_c_5 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 17 to port 5
R5_17 nt_n_17 nt_c_5 0.003124999999999963
X529 nt_n_17 nt_c_5 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X530 nt_p_17 nt_c_5 rl_admittance res=187800143092.54297 ind=8.409869753766284
X531 nt_p_17 nt_c_5 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X532 nt_p_17 nt_c_5 rl_admittance res=63732557064.23586 ind=35.261662271871394
X533 nt_n_17 nt_c_5 rl_admittance res=112799484372.98152 ind=31.919389834390056
X534 nt_n_17 nt_c_5 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 18 to port 5
R5_18 nt_n_18 nt_c_5 0.003124999999999963
X535 nt_n_18 nt_c_5 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X536 nt_p_18 nt_c_5 rl_admittance res=187800143092.54297 ind=8.409869753766284
X537 nt_p_18 nt_c_5 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X538 nt_p_18 nt_c_5 rl_admittance res=63732557064.23586 ind=35.261662271871394
X539 nt_n_18 nt_c_5 rl_admittance res=112799484372.98152 ind=31.919389834390056
X540 nt_n_18 nt_c_5 rl_admittance res=51262611157.92125 ind=93.72728905498322

* Port network for port 6
R_ref_6 p6 a6 50.0
H_b_6 a6 0 V_c_6 14.142135623730951
* Differential incident wave a sources for transfer from port 6
H_p_6 nt_p_6 nts_p_6 H_b_6 3.5355339059327378
E_p_6 nts_p_6 0 p6 0 0.07071067811865475
E_n_6 0 nt_n_6 nt_p_6 0 1
* Current sensor on center node for transfer to port 6
V_c_6 nt_c_6 0 0
* Transfer network from port 1 to port 6
R6_1 nt_n_1 nt_c_6 0.003124999999999963
X541 nt_n_1 nt_c_6 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X542 nt_p_1 nt_c_6 rl_admittance res=187800143092.54297 ind=8.409869753766284
X543 nt_p_1 nt_c_6 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X544 nt_p_1 nt_c_6 rl_admittance res=63732557064.23586 ind=35.261662271871394
X545 nt_n_1 nt_c_6 rl_admittance res=112799484372.98152 ind=31.919389834390056
X546 nt_n_1 nt_c_6 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 2 to port 6
R6_2 nt_n_2 nt_c_6 0.003124999999999963
X547 nt_n_2 nt_c_6 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X548 nt_p_2 nt_c_6 rl_admittance res=187800143092.54297 ind=8.409869753766284
X549 nt_p_2 nt_c_6 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X550 nt_p_2 nt_c_6 rl_admittance res=63732557064.23586 ind=35.261662271871394
X551 nt_n_2 nt_c_6 rl_admittance res=112799484372.98152 ind=31.919389834390056
X552 nt_n_2 nt_c_6 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 3 to port 6
R6_3 nt_n_3 nt_c_6 0.003124999999999963
X553 nt_n_3 nt_c_6 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X554 nt_p_3 nt_c_6 rl_admittance res=187800143092.54297 ind=8.409869753766284
X555 nt_p_3 nt_c_6 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X556 nt_p_3 nt_c_6 rl_admittance res=63732557064.23586 ind=35.261662271871394
X557 nt_n_3 nt_c_6 rl_admittance res=112799484372.98152 ind=31.919389834390056
X558 nt_n_3 nt_c_6 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 4 to port 6
R6_4 nt_n_4 nt_c_6 0.003124999999999963
X559 nt_n_4 nt_c_6 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X560 nt_p_4 nt_c_6 rl_admittance res=187800143092.54297 ind=8.409869753766284
X561 nt_p_4 nt_c_6 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X562 nt_p_4 nt_c_6 rl_admittance res=63732557064.23586 ind=35.261662271871394
X563 nt_n_4 nt_c_6 rl_admittance res=112799484372.98152 ind=31.919389834390056
X564 nt_n_4 nt_c_6 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 5 to port 6
R6_5 nt_n_5 nt_c_6 0.003124999999999963
X565 nt_n_5 nt_c_6 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X566 nt_p_5 nt_c_6 rl_admittance res=187800143092.54297 ind=8.409869753766284
X567 nt_p_5 nt_c_6 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X568 nt_p_5 nt_c_6 rl_admittance res=63732557064.23586 ind=35.261662271871394
X569 nt_n_5 nt_c_6 rl_admittance res=112799484372.98152 ind=31.919389834390056
X570 nt_n_5 nt_c_6 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 6 to port 6
R6_6 nt_p_6 nt_c_6 0.0007564900050830436
X571 nt_p_6 nt_c_6 rl_admittance res=6.713812060922877e+16 ind=0.01239433452121846
X572 nt_n_6 nt_c_6 rl_admittance res=0.00045787217518182793 ind=2.0503953265122565e-14
X573 nt_p_6 nt_c_6 rl_admittance res=0.00054254751817662 ind=7.679384261163742e-14
X574 nt_p_6 nt_c_6 rl_admittance res=0.0005564228350387422 ind=3.0785512135842906e-13
X575 nt_n_6 nt_c_6 rl_admittance res=0.0005055304090704312 ind=1.4305226916553906e-13
X576 nt_n_6 nt_c_6 rl_admittance res=0.00047272890640632993 ind=8.643258284073119e-13
* Transfer network from port 7 to port 6
R6_7 nt_n_7 nt_c_6 0.003124999999999963
X577 nt_n_7 nt_c_6 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X578 nt_p_7 nt_c_6 rl_admittance res=187800143092.54297 ind=8.409869753766284
X579 nt_p_7 nt_c_6 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X580 nt_p_7 nt_c_6 rl_admittance res=63732557064.23586 ind=35.261662271871394
X581 nt_n_7 nt_c_6 rl_admittance res=112799484372.98152 ind=31.919389834390056
X582 nt_n_7 nt_c_6 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 8 to port 6
R6_8 nt_n_8 nt_c_6 0.003124999999999963
X583 nt_n_8 nt_c_6 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X584 nt_p_8 nt_c_6 rl_admittance res=187800143092.54297 ind=8.409869753766284
X585 nt_p_8 nt_c_6 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X586 nt_p_8 nt_c_6 rl_admittance res=63732557064.23586 ind=35.261662271871394
X587 nt_n_8 nt_c_6 rl_admittance res=112799484372.98152 ind=31.919389834390056
X588 nt_n_8 nt_c_6 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 9 to port 6
R6_9 nt_n_9 nt_c_6 0.003124999999999963
X589 nt_n_9 nt_c_6 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X590 nt_p_9 nt_c_6 rl_admittance res=187800143092.54297 ind=8.409869753766284
X591 nt_p_9 nt_c_6 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X592 nt_p_9 nt_c_6 rl_admittance res=63732557064.23586 ind=35.261662271871394
X593 nt_n_9 nt_c_6 rl_admittance res=112799484372.98152 ind=31.919389834390056
X594 nt_n_9 nt_c_6 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 10 to port 6
R6_10 nt_n_10 nt_c_6 0.003124999999999963
X595 nt_n_10 nt_c_6 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X596 nt_p_10 nt_c_6 rl_admittance res=187800143092.54297 ind=8.409869753766284
X597 nt_p_10 nt_c_6 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X598 nt_p_10 nt_c_6 rl_admittance res=63732557064.23586 ind=35.261662271871394
X599 nt_n_10 nt_c_6 rl_admittance res=112799484372.98152 ind=31.919389834390056
X600 nt_n_10 nt_c_6 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 11 to port 6
R6_11 nt_n_11 nt_c_6 0.003124999999999963
X601 nt_n_11 nt_c_6 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X602 nt_p_11 nt_c_6 rl_admittance res=187800143092.54297 ind=8.409869753766284
X603 nt_p_11 nt_c_6 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X604 nt_p_11 nt_c_6 rl_admittance res=63732557064.23586 ind=35.261662271871394
X605 nt_n_11 nt_c_6 rl_admittance res=112799484372.98152 ind=31.919389834390056
X606 nt_n_11 nt_c_6 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 12 to port 6
R6_12 nt_n_12 nt_c_6 0.003124999999999963
X607 nt_n_12 nt_c_6 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X608 nt_p_12 nt_c_6 rl_admittance res=187800143092.54297 ind=8.409869753766284
X609 nt_p_12 nt_c_6 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X610 nt_p_12 nt_c_6 rl_admittance res=63732557064.23586 ind=35.261662271871394
X611 nt_n_12 nt_c_6 rl_admittance res=112799484372.98152 ind=31.919389834390056
X612 nt_n_12 nt_c_6 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 13 to port 6
R6_13 nt_n_13 nt_c_6 0.003124999999999963
X613 nt_n_13 nt_c_6 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X614 nt_p_13 nt_c_6 rl_admittance res=187800143092.54297 ind=8.409869753766284
X615 nt_p_13 nt_c_6 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X616 nt_p_13 nt_c_6 rl_admittance res=63732557064.23586 ind=35.261662271871394
X617 nt_n_13 nt_c_6 rl_admittance res=112799484372.98152 ind=31.919389834390056
X618 nt_n_13 nt_c_6 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 14 to port 6
R6_14 nt_n_14 nt_c_6 0.003124999999999963
X619 nt_n_14 nt_c_6 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X620 nt_p_14 nt_c_6 rl_admittance res=187800143092.54297 ind=8.409869753766284
X621 nt_p_14 nt_c_6 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X622 nt_p_14 nt_c_6 rl_admittance res=63732557064.23586 ind=35.261662271871394
X623 nt_n_14 nt_c_6 rl_admittance res=112799484372.98152 ind=31.919389834390056
X624 nt_n_14 nt_c_6 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 15 to port 6
R6_15 nt_n_15 nt_c_6 0.003124999999999963
X625 nt_n_15 nt_c_6 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X626 nt_p_15 nt_c_6 rl_admittance res=187800143092.54297 ind=8.409869753766284
X627 nt_p_15 nt_c_6 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X628 nt_p_15 nt_c_6 rl_admittance res=63732557064.23586 ind=35.261662271871394
X629 nt_n_15 nt_c_6 rl_admittance res=112799484372.98152 ind=31.919389834390056
X630 nt_n_15 nt_c_6 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 16 to port 6
R6_16 nt_n_16 nt_c_6 0.003124999999999963
X631 nt_n_16 nt_c_6 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X632 nt_p_16 nt_c_6 rl_admittance res=187800143092.54297 ind=8.409869753766284
X633 nt_p_16 nt_c_6 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X634 nt_p_16 nt_c_6 rl_admittance res=63732557064.23586 ind=35.261662271871394
X635 nt_n_16 nt_c_6 rl_admittance res=112799484372.98152 ind=31.919389834390056
X636 nt_n_16 nt_c_6 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 17 to port 6
R6_17 nt_n_17 nt_c_6 0.003124999999999963
X637 nt_n_17 nt_c_6 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X638 nt_p_17 nt_c_6 rl_admittance res=187800143092.54297 ind=8.409869753766284
X639 nt_p_17 nt_c_6 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X640 nt_p_17 nt_c_6 rl_admittance res=63732557064.23586 ind=35.261662271871394
X641 nt_n_17 nt_c_6 rl_admittance res=112799484372.98152 ind=31.919389834390056
X642 nt_n_17 nt_c_6 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 18 to port 6
R6_18 nt_n_18 nt_c_6 0.003124999999999963
X643 nt_n_18 nt_c_6 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X644 nt_p_18 nt_c_6 rl_admittance res=187800143092.54297 ind=8.409869753766284
X645 nt_p_18 nt_c_6 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X646 nt_p_18 nt_c_6 rl_admittance res=63732557064.23586 ind=35.261662271871394
X647 nt_n_18 nt_c_6 rl_admittance res=112799484372.98152 ind=31.919389834390056
X648 nt_n_18 nt_c_6 rl_admittance res=51262611157.92125 ind=93.72728905498322

* Port network for port 7
R_ref_7 p7 a7 50.0
H_b_7 a7 0 V_c_7 14.142135623730951
* Differential incident wave a sources for transfer from port 7
H_p_7 nt_p_7 nts_p_7 H_b_7 3.5355339059327378
E_p_7 nts_p_7 0 p7 0 0.07071067811865475
E_n_7 0 nt_n_7 nt_p_7 0 1
* Current sensor on center node for transfer to port 7
V_c_7 nt_c_7 0 0
* Transfer network from port 1 to port 7
R7_1 nt_n_1 nt_c_7 0.003124999999999963
X649 nt_n_1 nt_c_7 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X650 nt_p_1 nt_c_7 rl_admittance res=187800143092.54297 ind=8.409869753766284
X651 nt_p_1 nt_c_7 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X652 nt_p_1 nt_c_7 rl_admittance res=63732557064.23586 ind=35.261662271871394
X653 nt_n_1 nt_c_7 rl_admittance res=112799484372.98152 ind=31.919389834390056
X654 nt_n_1 nt_c_7 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 2 to port 7
R7_2 nt_n_2 nt_c_7 0.003124999999999963
X655 nt_n_2 nt_c_7 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X656 nt_p_2 nt_c_7 rl_admittance res=187800143092.54297 ind=8.409869753766284
X657 nt_p_2 nt_c_7 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X658 nt_p_2 nt_c_7 rl_admittance res=63732557064.23586 ind=35.261662271871394
X659 nt_n_2 nt_c_7 rl_admittance res=112799484372.98152 ind=31.919389834390056
X660 nt_n_2 nt_c_7 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 3 to port 7
R7_3 nt_n_3 nt_c_7 0.003124999999999963
X661 nt_n_3 nt_c_7 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X662 nt_p_3 nt_c_7 rl_admittance res=187800143092.54297 ind=8.409869753766284
X663 nt_p_3 nt_c_7 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X664 nt_p_3 nt_c_7 rl_admittance res=63732557064.23586 ind=35.261662271871394
X665 nt_n_3 nt_c_7 rl_admittance res=112799484372.98152 ind=31.919389834390056
X666 nt_n_3 nt_c_7 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 4 to port 7
R7_4 nt_n_4 nt_c_7 0.003124999999999963
X667 nt_n_4 nt_c_7 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X668 nt_p_4 nt_c_7 rl_admittance res=187800143092.54297 ind=8.409869753766284
X669 nt_p_4 nt_c_7 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X670 nt_p_4 nt_c_7 rl_admittance res=63732557064.23586 ind=35.261662271871394
X671 nt_n_4 nt_c_7 rl_admittance res=112799484372.98152 ind=31.919389834390056
X672 nt_n_4 nt_c_7 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 5 to port 7
R7_5 nt_n_5 nt_c_7 0.003124999999999963
X673 nt_n_5 nt_c_7 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X674 nt_p_5 nt_c_7 rl_admittance res=187800143092.54297 ind=8.409869753766284
X675 nt_p_5 nt_c_7 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X676 nt_p_5 nt_c_7 rl_admittance res=63732557064.23586 ind=35.261662271871394
X677 nt_n_5 nt_c_7 rl_admittance res=112799484372.98152 ind=31.919389834390056
X678 nt_n_5 nt_c_7 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 6 to port 7
R7_6 nt_n_6 nt_c_7 0.003124999999999963
X679 nt_n_6 nt_c_7 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X680 nt_p_6 nt_c_7 rl_admittance res=187800143092.54297 ind=8.409869753766284
X681 nt_p_6 nt_c_7 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X682 nt_p_6 nt_c_7 rl_admittance res=63732557064.23586 ind=35.261662271871394
X683 nt_n_6 nt_c_7 rl_admittance res=112799484372.98152 ind=31.919389834390056
X684 nt_n_6 nt_c_7 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 7 to port 7
R7_7 nt_p_7 nt_c_7 0.0007564900050830436
X685 nt_p_7 nt_c_7 rl_admittance res=6.713812060922877e+16 ind=0.01239433452121846
X686 nt_n_7 nt_c_7 rl_admittance res=0.00045787217518182793 ind=2.0503953265122565e-14
X687 nt_p_7 nt_c_7 rl_admittance res=0.00054254751817662 ind=7.679384261163742e-14
X688 nt_p_7 nt_c_7 rl_admittance res=0.0005564228350387422 ind=3.0785512135842906e-13
X689 nt_n_7 nt_c_7 rl_admittance res=0.0005055304090704312 ind=1.4305226916553906e-13
X690 nt_n_7 nt_c_7 rl_admittance res=0.00047272890640632993 ind=8.643258284073119e-13
* Transfer network from port 8 to port 7
R7_8 nt_n_8 nt_c_7 0.003124999999999963
X691 nt_n_8 nt_c_7 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X692 nt_p_8 nt_c_7 rl_admittance res=187800143092.54297 ind=8.409869753766284
X693 nt_p_8 nt_c_7 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X694 nt_p_8 nt_c_7 rl_admittance res=63732557064.23586 ind=35.261662271871394
X695 nt_n_8 nt_c_7 rl_admittance res=112799484372.98152 ind=31.919389834390056
X696 nt_n_8 nt_c_7 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 9 to port 7
R7_9 nt_n_9 nt_c_7 0.003124999999999963
X697 nt_n_9 nt_c_7 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X698 nt_p_9 nt_c_7 rl_admittance res=187800143092.54297 ind=8.409869753766284
X699 nt_p_9 nt_c_7 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X700 nt_p_9 nt_c_7 rl_admittance res=63732557064.23586 ind=35.261662271871394
X701 nt_n_9 nt_c_7 rl_admittance res=112799484372.98152 ind=31.919389834390056
X702 nt_n_9 nt_c_7 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 10 to port 7
R7_10 nt_n_10 nt_c_7 0.003124999999999963
X703 nt_n_10 nt_c_7 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X704 nt_p_10 nt_c_7 rl_admittance res=187800143092.54297 ind=8.409869753766284
X705 nt_p_10 nt_c_7 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X706 nt_p_10 nt_c_7 rl_admittance res=63732557064.23586 ind=35.261662271871394
X707 nt_n_10 nt_c_7 rl_admittance res=112799484372.98152 ind=31.919389834390056
X708 nt_n_10 nt_c_7 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 11 to port 7
R7_11 nt_n_11 nt_c_7 0.003124999999999963
X709 nt_n_11 nt_c_7 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X710 nt_p_11 nt_c_7 rl_admittance res=187800143092.54297 ind=8.409869753766284
X711 nt_p_11 nt_c_7 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X712 nt_p_11 nt_c_7 rl_admittance res=63732557064.23586 ind=35.261662271871394
X713 nt_n_11 nt_c_7 rl_admittance res=112799484372.98152 ind=31.919389834390056
X714 nt_n_11 nt_c_7 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 12 to port 7
R7_12 nt_n_12 nt_c_7 0.003124999999999963
X715 nt_n_12 nt_c_7 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X716 nt_p_12 nt_c_7 rl_admittance res=187800143092.54297 ind=8.409869753766284
X717 nt_p_12 nt_c_7 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X718 nt_p_12 nt_c_7 rl_admittance res=63732557064.23586 ind=35.261662271871394
X719 nt_n_12 nt_c_7 rl_admittance res=112799484372.98152 ind=31.919389834390056
X720 nt_n_12 nt_c_7 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 13 to port 7
R7_13 nt_n_13 nt_c_7 0.003124999999999963
X721 nt_n_13 nt_c_7 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X722 nt_p_13 nt_c_7 rl_admittance res=187800143092.54297 ind=8.409869753766284
X723 nt_p_13 nt_c_7 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X724 nt_p_13 nt_c_7 rl_admittance res=63732557064.23586 ind=35.261662271871394
X725 nt_n_13 nt_c_7 rl_admittance res=112799484372.98152 ind=31.919389834390056
X726 nt_n_13 nt_c_7 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 14 to port 7
R7_14 nt_n_14 nt_c_7 0.003124999999999963
X727 nt_n_14 nt_c_7 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X728 nt_p_14 nt_c_7 rl_admittance res=187800143092.54297 ind=8.409869753766284
X729 nt_p_14 nt_c_7 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X730 nt_p_14 nt_c_7 rl_admittance res=63732557064.23586 ind=35.261662271871394
X731 nt_n_14 nt_c_7 rl_admittance res=112799484372.98152 ind=31.919389834390056
X732 nt_n_14 nt_c_7 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 15 to port 7
R7_15 nt_n_15 nt_c_7 0.003124999999999963
X733 nt_n_15 nt_c_7 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X734 nt_p_15 nt_c_7 rl_admittance res=187800143092.54297 ind=8.409869753766284
X735 nt_p_15 nt_c_7 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X736 nt_p_15 nt_c_7 rl_admittance res=63732557064.23586 ind=35.261662271871394
X737 nt_n_15 nt_c_7 rl_admittance res=112799484372.98152 ind=31.919389834390056
X738 nt_n_15 nt_c_7 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 16 to port 7
R7_16 nt_n_16 nt_c_7 0.003124999999999963
X739 nt_n_16 nt_c_7 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X740 nt_p_16 nt_c_7 rl_admittance res=187800143092.54297 ind=8.409869753766284
X741 nt_p_16 nt_c_7 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X742 nt_p_16 nt_c_7 rl_admittance res=63732557064.23586 ind=35.261662271871394
X743 nt_n_16 nt_c_7 rl_admittance res=112799484372.98152 ind=31.919389834390056
X744 nt_n_16 nt_c_7 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 17 to port 7
R7_17 nt_n_17 nt_c_7 0.003124999999999963
X745 nt_n_17 nt_c_7 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X746 nt_p_17 nt_c_7 rl_admittance res=187800143092.54297 ind=8.409869753766284
X747 nt_p_17 nt_c_7 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X748 nt_p_17 nt_c_7 rl_admittance res=63732557064.23586 ind=35.261662271871394
X749 nt_n_17 nt_c_7 rl_admittance res=112799484372.98152 ind=31.919389834390056
X750 nt_n_17 nt_c_7 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 18 to port 7
R7_18 nt_n_18 nt_c_7 0.003124999999999963
X751 nt_n_18 nt_c_7 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X752 nt_p_18 nt_c_7 rl_admittance res=187800143092.54297 ind=8.409869753766284
X753 nt_p_18 nt_c_7 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X754 nt_p_18 nt_c_7 rl_admittance res=63732557064.23586 ind=35.261662271871394
X755 nt_n_18 nt_c_7 rl_admittance res=112799484372.98152 ind=31.919389834390056
X756 nt_n_18 nt_c_7 rl_admittance res=51262611157.92125 ind=93.72728905498322

* Port network for port 8
R_ref_8 p8 a8 50.0
H_b_8 a8 0 V_c_8 14.142135623730951
* Differential incident wave a sources for transfer from port 8
H_p_8 nt_p_8 nts_p_8 H_b_8 3.5355339059327378
E_p_8 nts_p_8 0 p8 0 0.07071067811865475
E_n_8 0 nt_n_8 nt_p_8 0 1
* Current sensor on center node for transfer to port 8
V_c_8 nt_c_8 0 0
* Transfer network from port 1 to port 8
R8_1 nt_n_1 nt_c_8 0.003124999999999963
X757 nt_n_1 nt_c_8 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X758 nt_p_1 nt_c_8 rl_admittance res=187800143092.54297 ind=8.409869753766284
X759 nt_p_1 nt_c_8 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X760 nt_p_1 nt_c_8 rl_admittance res=63732557064.23586 ind=35.261662271871394
X761 nt_n_1 nt_c_8 rl_admittance res=112799484372.98152 ind=31.919389834390056
X762 nt_n_1 nt_c_8 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 2 to port 8
R8_2 nt_n_2 nt_c_8 0.003124999999999963
X763 nt_n_2 nt_c_8 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X764 nt_p_2 nt_c_8 rl_admittance res=187800143092.54297 ind=8.409869753766284
X765 nt_p_2 nt_c_8 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X766 nt_p_2 nt_c_8 rl_admittance res=63732557064.23586 ind=35.261662271871394
X767 nt_n_2 nt_c_8 rl_admittance res=112799484372.98152 ind=31.919389834390056
X768 nt_n_2 nt_c_8 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 3 to port 8
R8_3 nt_n_3 nt_c_8 0.003124999999999963
X769 nt_n_3 nt_c_8 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X770 nt_p_3 nt_c_8 rl_admittance res=187800143092.54297 ind=8.409869753766284
X771 nt_p_3 nt_c_8 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X772 nt_p_3 nt_c_8 rl_admittance res=63732557064.23586 ind=35.261662271871394
X773 nt_n_3 nt_c_8 rl_admittance res=112799484372.98152 ind=31.919389834390056
X774 nt_n_3 nt_c_8 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 4 to port 8
R8_4 nt_n_4 nt_c_8 0.003124999999999963
X775 nt_n_4 nt_c_8 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X776 nt_p_4 nt_c_8 rl_admittance res=187800143092.54297 ind=8.409869753766284
X777 nt_p_4 nt_c_8 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X778 nt_p_4 nt_c_8 rl_admittance res=63732557064.23586 ind=35.261662271871394
X779 nt_n_4 nt_c_8 rl_admittance res=112799484372.98152 ind=31.919389834390056
X780 nt_n_4 nt_c_8 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 5 to port 8
R8_5 nt_n_5 nt_c_8 0.003124999999999963
X781 nt_n_5 nt_c_8 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X782 nt_p_5 nt_c_8 rl_admittance res=187800143092.54297 ind=8.409869753766284
X783 nt_p_5 nt_c_8 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X784 nt_p_5 nt_c_8 rl_admittance res=63732557064.23586 ind=35.261662271871394
X785 nt_n_5 nt_c_8 rl_admittance res=112799484372.98152 ind=31.919389834390056
X786 nt_n_5 nt_c_8 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 6 to port 8
R8_6 nt_n_6 nt_c_8 0.003124999999999963
X787 nt_n_6 nt_c_8 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X788 nt_p_6 nt_c_8 rl_admittance res=187800143092.54297 ind=8.409869753766284
X789 nt_p_6 nt_c_8 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X790 nt_p_6 nt_c_8 rl_admittance res=63732557064.23586 ind=35.261662271871394
X791 nt_n_6 nt_c_8 rl_admittance res=112799484372.98152 ind=31.919389834390056
X792 nt_n_6 nt_c_8 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 7 to port 8
R8_7 nt_n_7 nt_c_8 0.003124999999999963
X793 nt_n_7 nt_c_8 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X794 nt_p_7 nt_c_8 rl_admittance res=187800143092.54297 ind=8.409869753766284
X795 nt_p_7 nt_c_8 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X796 nt_p_7 nt_c_8 rl_admittance res=63732557064.23586 ind=35.261662271871394
X797 nt_n_7 nt_c_8 rl_admittance res=112799484372.98152 ind=31.919389834390056
X798 nt_n_7 nt_c_8 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 8 to port 8
R8_8 nt_p_8 nt_c_8 0.0007564900050830436
X799 nt_p_8 nt_c_8 rl_admittance res=6.713812060922877e+16 ind=0.01239433452121846
X800 nt_n_8 nt_c_8 rl_admittance res=0.00045787217518182793 ind=2.0503953265122565e-14
X801 nt_p_8 nt_c_8 rl_admittance res=0.00054254751817662 ind=7.679384261163742e-14
X802 nt_p_8 nt_c_8 rl_admittance res=0.0005564228350387422 ind=3.0785512135842906e-13
X803 nt_n_8 nt_c_8 rl_admittance res=0.0005055304090704312 ind=1.4305226916553906e-13
X804 nt_n_8 nt_c_8 rl_admittance res=0.00047272890640632993 ind=8.643258284073119e-13
* Transfer network from port 9 to port 8
R8_9 nt_n_9 nt_c_8 0.003124999999999963
X805 nt_n_9 nt_c_8 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X806 nt_p_9 nt_c_8 rl_admittance res=187800143092.54297 ind=8.409869753766284
X807 nt_p_9 nt_c_8 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X808 nt_p_9 nt_c_8 rl_admittance res=63732557064.23586 ind=35.261662271871394
X809 nt_n_9 nt_c_8 rl_admittance res=112799484372.98152 ind=31.919389834390056
X810 nt_n_9 nt_c_8 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 10 to port 8
R8_10 nt_n_10 nt_c_8 0.003124999999999963
X811 nt_n_10 nt_c_8 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X812 nt_p_10 nt_c_8 rl_admittance res=187800143092.54297 ind=8.409869753766284
X813 nt_p_10 nt_c_8 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X814 nt_p_10 nt_c_8 rl_admittance res=63732557064.23586 ind=35.261662271871394
X815 nt_n_10 nt_c_8 rl_admittance res=112799484372.98152 ind=31.919389834390056
X816 nt_n_10 nt_c_8 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 11 to port 8
R8_11 nt_n_11 nt_c_8 0.003124999999999963
X817 nt_n_11 nt_c_8 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X818 nt_p_11 nt_c_8 rl_admittance res=187800143092.54297 ind=8.409869753766284
X819 nt_p_11 nt_c_8 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X820 nt_p_11 nt_c_8 rl_admittance res=63732557064.23586 ind=35.261662271871394
X821 nt_n_11 nt_c_8 rl_admittance res=112799484372.98152 ind=31.919389834390056
X822 nt_n_11 nt_c_8 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 12 to port 8
R8_12 nt_n_12 nt_c_8 0.003124999999999963
X823 nt_n_12 nt_c_8 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X824 nt_p_12 nt_c_8 rl_admittance res=187800143092.54297 ind=8.409869753766284
X825 nt_p_12 nt_c_8 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X826 nt_p_12 nt_c_8 rl_admittance res=63732557064.23586 ind=35.261662271871394
X827 nt_n_12 nt_c_8 rl_admittance res=112799484372.98152 ind=31.919389834390056
X828 nt_n_12 nt_c_8 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 13 to port 8
R8_13 nt_n_13 nt_c_8 0.003124999999999963
X829 nt_n_13 nt_c_8 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X830 nt_p_13 nt_c_8 rl_admittance res=187800143092.54297 ind=8.409869753766284
X831 nt_p_13 nt_c_8 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X832 nt_p_13 nt_c_8 rl_admittance res=63732557064.23586 ind=35.261662271871394
X833 nt_n_13 nt_c_8 rl_admittance res=112799484372.98152 ind=31.919389834390056
X834 nt_n_13 nt_c_8 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 14 to port 8
R8_14 nt_n_14 nt_c_8 0.003124999999999963
X835 nt_n_14 nt_c_8 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X836 nt_p_14 nt_c_8 rl_admittance res=187800143092.54297 ind=8.409869753766284
X837 nt_p_14 nt_c_8 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X838 nt_p_14 nt_c_8 rl_admittance res=63732557064.23586 ind=35.261662271871394
X839 nt_n_14 nt_c_8 rl_admittance res=112799484372.98152 ind=31.919389834390056
X840 nt_n_14 nt_c_8 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 15 to port 8
R8_15 nt_n_15 nt_c_8 0.003124999999999963
X841 nt_n_15 nt_c_8 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X842 nt_p_15 nt_c_8 rl_admittance res=187800143092.54297 ind=8.409869753766284
X843 nt_p_15 nt_c_8 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X844 nt_p_15 nt_c_8 rl_admittance res=63732557064.23586 ind=35.261662271871394
X845 nt_n_15 nt_c_8 rl_admittance res=112799484372.98152 ind=31.919389834390056
X846 nt_n_15 nt_c_8 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 16 to port 8
R8_16 nt_n_16 nt_c_8 0.003124999999999963
X847 nt_n_16 nt_c_8 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X848 nt_p_16 nt_c_8 rl_admittance res=187800143092.54297 ind=8.409869753766284
X849 nt_p_16 nt_c_8 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X850 nt_p_16 nt_c_8 rl_admittance res=63732557064.23586 ind=35.261662271871394
X851 nt_n_16 nt_c_8 rl_admittance res=112799484372.98152 ind=31.919389834390056
X852 nt_n_16 nt_c_8 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 17 to port 8
R8_17 nt_n_17 nt_c_8 0.003124999999999963
X853 nt_n_17 nt_c_8 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X854 nt_p_17 nt_c_8 rl_admittance res=187800143092.54297 ind=8.409869753766284
X855 nt_p_17 nt_c_8 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X856 nt_p_17 nt_c_8 rl_admittance res=63732557064.23586 ind=35.261662271871394
X857 nt_n_17 nt_c_8 rl_admittance res=112799484372.98152 ind=31.919389834390056
X858 nt_n_17 nt_c_8 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 18 to port 8
R8_18 nt_n_18 nt_c_8 0.003124999999999963
X859 nt_n_18 nt_c_8 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X860 nt_p_18 nt_c_8 rl_admittance res=187800143092.54297 ind=8.409869753766284
X861 nt_p_18 nt_c_8 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X862 nt_p_18 nt_c_8 rl_admittance res=63732557064.23586 ind=35.261662271871394
X863 nt_n_18 nt_c_8 rl_admittance res=112799484372.98152 ind=31.919389834390056
X864 nt_n_18 nt_c_8 rl_admittance res=51262611157.92125 ind=93.72728905498322

* Port network for port 9
R_ref_9 p9 a9 50.0
H_b_9 a9 0 V_c_9 14.142135623730951
* Differential incident wave a sources for transfer from port 9
H_p_9 nt_p_9 nts_p_9 H_b_9 3.5355339059327378
E_p_9 nts_p_9 0 p9 0 0.07071067811865475
E_n_9 0 nt_n_9 nt_p_9 0 1
* Current sensor on center node for transfer to port 9
V_c_9 nt_c_9 0 0
* Transfer network from port 1 to port 9
R9_1 nt_n_1 nt_c_9 0.003124999999999963
X865 nt_n_1 nt_c_9 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X866 nt_p_1 nt_c_9 rl_admittance res=187800143092.54297 ind=8.409869753766284
X867 nt_p_1 nt_c_9 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X868 nt_p_1 nt_c_9 rl_admittance res=63732557064.23586 ind=35.261662271871394
X869 nt_n_1 nt_c_9 rl_admittance res=112799484372.98152 ind=31.919389834390056
X870 nt_n_1 nt_c_9 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 2 to port 9
R9_2 nt_n_2 nt_c_9 0.003124999999999963
X871 nt_n_2 nt_c_9 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X872 nt_p_2 nt_c_9 rl_admittance res=187800143092.54297 ind=8.409869753766284
X873 nt_p_2 nt_c_9 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X874 nt_p_2 nt_c_9 rl_admittance res=63732557064.23586 ind=35.261662271871394
X875 nt_n_2 nt_c_9 rl_admittance res=112799484372.98152 ind=31.919389834390056
X876 nt_n_2 nt_c_9 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 3 to port 9
R9_3 nt_n_3 nt_c_9 0.003124999999999963
X877 nt_n_3 nt_c_9 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X878 nt_p_3 nt_c_9 rl_admittance res=187800143092.54297 ind=8.409869753766284
X879 nt_p_3 nt_c_9 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X880 nt_p_3 nt_c_9 rl_admittance res=63732557064.23586 ind=35.261662271871394
X881 nt_n_3 nt_c_9 rl_admittance res=112799484372.98152 ind=31.919389834390056
X882 nt_n_3 nt_c_9 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 4 to port 9
R9_4 nt_n_4 nt_c_9 0.003124999999999963
X883 nt_n_4 nt_c_9 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X884 nt_p_4 nt_c_9 rl_admittance res=187800143092.54297 ind=8.409869753766284
X885 nt_p_4 nt_c_9 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X886 nt_p_4 nt_c_9 rl_admittance res=63732557064.23586 ind=35.261662271871394
X887 nt_n_4 nt_c_9 rl_admittance res=112799484372.98152 ind=31.919389834390056
X888 nt_n_4 nt_c_9 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 5 to port 9
R9_5 nt_n_5 nt_c_9 0.003124999999999963
X889 nt_n_5 nt_c_9 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X890 nt_p_5 nt_c_9 rl_admittance res=187800143092.54297 ind=8.409869753766284
X891 nt_p_5 nt_c_9 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X892 nt_p_5 nt_c_9 rl_admittance res=63732557064.23586 ind=35.261662271871394
X893 nt_n_5 nt_c_9 rl_admittance res=112799484372.98152 ind=31.919389834390056
X894 nt_n_5 nt_c_9 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 6 to port 9
R9_6 nt_n_6 nt_c_9 0.003124999999999963
X895 nt_n_6 nt_c_9 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X896 nt_p_6 nt_c_9 rl_admittance res=187800143092.54297 ind=8.409869753766284
X897 nt_p_6 nt_c_9 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X898 nt_p_6 nt_c_9 rl_admittance res=63732557064.23586 ind=35.261662271871394
X899 nt_n_6 nt_c_9 rl_admittance res=112799484372.98152 ind=31.919389834390056
X900 nt_n_6 nt_c_9 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 7 to port 9
R9_7 nt_n_7 nt_c_9 0.003124999999999963
X901 nt_n_7 nt_c_9 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X902 nt_p_7 nt_c_9 rl_admittance res=187800143092.54297 ind=8.409869753766284
X903 nt_p_7 nt_c_9 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X904 nt_p_7 nt_c_9 rl_admittance res=63732557064.23586 ind=35.261662271871394
X905 nt_n_7 nt_c_9 rl_admittance res=112799484372.98152 ind=31.919389834390056
X906 nt_n_7 nt_c_9 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 8 to port 9
R9_8 nt_n_8 nt_c_9 0.003124999999999963
X907 nt_n_8 nt_c_9 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X908 nt_p_8 nt_c_9 rl_admittance res=187800143092.54297 ind=8.409869753766284
X909 nt_p_8 nt_c_9 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X910 nt_p_8 nt_c_9 rl_admittance res=63732557064.23586 ind=35.261662271871394
X911 nt_n_8 nt_c_9 rl_admittance res=112799484372.98152 ind=31.919389834390056
X912 nt_n_8 nt_c_9 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 9 to port 9
R9_9 nt_p_9 nt_c_9 0.0007564900050830436
X913 nt_p_9 nt_c_9 rl_admittance res=6.713812060922877e+16 ind=0.01239433452121846
X914 nt_n_9 nt_c_9 rl_admittance res=0.00045787217518182793 ind=2.0503953265122565e-14
X915 nt_p_9 nt_c_9 rl_admittance res=0.00054254751817662 ind=7.679384261163742e-14
X916 nt_p_9 nt_c_9 rl_admittance res=0.0005564228350387422 ind=3.0785512135842906e-13
X917 nt_n_9 nt_c_9 rl_admittance res=0.0005055304090704312 ind=1.4305226916553906e-13
X918 nt_n_9 nt_c_9 rl_admittance res=0.00047272890640632993 ind=8.643258284073119e-13
* Transfer network from port 10 to port 9
R9_10 nt_n_10 nt_c_9 0.003124999999999963
X919 nt_n_10 nt_c_9 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X920 nt_p_10 nt_c_9 rl_admittance res=187800143092.54297 ind=8.409869753766284
X921 nt_p_10 nt_c_9 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X922 nt_p_10 nt_c_9 rl_admittance res=63732557064.23586 ind=35.261662271871394
X923 nt_n_10 nt_c_9 rl_admittance res=112799484372.98152 ind=31.919389834390056
X924 nt_n_10 nt_c_9 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 11 to port 9
R9_11 nt_n_11 nt_c_9 0.003124999999999963
X925 nt_n_11 nt_c_9 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X926 nt_p_11 nt_c_9 rl_admittance res=187800143092.54297 ind=8.409869753766284
X927 nt_p_11 nt_c_9 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X928 nt_p_11 nt_c_9 rl_admittance res=63732557064.23586 ind=35.261662271871394
X929 nt_n_11 nt_c_9 rl_admittance res=112799484372.98152 ind=31.919389834390056
X930 nt_n_11 nt_c_9 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 12 to port 9
R9_12 nt_n_12 nt_c_9 0.003124999999999963
X931 nt_n_12 nt_c_9 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X932 nt_p_12 nt_c_9 rl_admittance res=187800143092.54297 ind=8.409869753766284
X933 nt_p_12 nt_c_9 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X934 nt_p_12 nt_c_9 rl_admittance res=63732557064.23586 ind=35.261662271871394
X935 nt_n_12 nt_c_9 rl_admittance res=112799484372.98152 ind=31.919389834390056
X936 nt_n_12 nt_c_9 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 13 to port 9
R9_13 nt_n_13 nt_c_9 0.003124999999999963
X937 nt_n_13 nt_c_9 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X938 nt_p_13 nt_c_9 rl_admittance res=187800143092.54297 ind=8.409869753766284
X939 nt_p_13 nt_c_9 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X940 nt_p_13 nt_c_9 rl_admittance res=63732557064.23586 ind=35.261662271871394
X941 nt_n_13 nt_c_9 rl_admittance res=112799484372.98152 ind=31.919389834390056
X942 nt_n_13 nt_c_9 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 14 to port 9
R9_14 nt_n_14 nt_c_9 0.003124999999999963
X943 nt_n_14 nt_c_9 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X944 nt_p_14 nt_c_9 rl_admittance res=187800143092.54297 ind=8.409869753766284
X945 nt_p_14 nt_c_9 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X946 nt_p_14 nt_c_9 rl_admittance res=63732557064.23586 ind=35.261662271871394
X947 nt_n_14 nt_c_9 rl_admittance res=112799484372.98152 ind=31.919389834390056
X948 nt_n_14 nt_c_9 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 15 to port 9
R9_15 nt_n_15 nt_c_9 0.003124999999999963
X949 nt_n_15 nt_c_9 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X950 nt_p_15 nt_c_9 rl_admittance res=187800143092.54297 ind=8.409869753766284
X951 nt_p_15 nt_c_9 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X952 nt_p_15 nt_c_9 rl_admittance res=63732557064.23586 ind=35.261662271871394
X953 nt_n_15 nt_c_9 rl_admittance res=112799484372.98152 ind=31.919389834390056
X954 nt_n_15 nt_c_9 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 16 to port 9
R9_16 nt_n_16 nt_c_9 0.003124999999999963
X955 nt_n_16 nt_c_9 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X956 nt_p_16 nt_c_9 rl_admittance res=187800143092.54297 ind=8.409869753766284
X957 nt_p_16 nt_c_9 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X958 nt_p_16 nt_c_9 rl_admittance res=63732557064.23586 ind=35.261662271871394
X959 nt_n_16 nt_c_9 rl_admittance res=112799484372.98152 ind=31.919389834390056
X960 nt_n_16 nt_c_9 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 17 to port 9
R9_17 nt_n_17 nt_c_9 0.003124999999999963
X961 nt_n_17 nt_c_9 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X962 nt_p_17 nt_c_9 rl_admittance res=187800143092.54297 ind=8.409869753766284
X963 nt_p_17 nt_c_9 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X964 nt_p_17 nt_c_9 rl_admittance res=63732557064.23586 ind=35.261662271871394
X965 nt_n_17 nt_c_9 rl_admittance res=112799484372.98152 ind=31.919389834390056
X966 nt_n_17 nt_c_9 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 18 to port 9
R9_18 nt_n_18 nt_c_9 0.003124999999999963
X967 nt_n_18 nt_c_9 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X968 nt_p_18 nt_c_9 rl_admittance res=187800143092.54297 ind=8.409869753766284
X969 nt_p_18 nt_c_9 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X970 nt_p_18 nt_c_9 rl_admittance res=63732557064.23586 ind=35.261662271871394
X971 nt_n_18 nt_c_9 rl_admittance res=112799484372.98152 ind=31.919389834390056
X972 nt_n_18 nt_c_9 rl_admittance res=51262611157.92125 ind=93.72728905498322

* Port network for port 10
R_ref_10 p10 a10 50.0
H_b_10 a10 0 V_c_10 14.142135623730951
* Differential incident wave a sources for transfer from port 10
H_p_10 nt_p_10 nts_p_10 H_b_10 3.5355339059327378
E_p_10 nts_p_10 0 p10 0 0.07071067811865475
E_n_10 0 nt_n_10 nt_p_10 0 1
* Current sensor on center node for transfer to port 10
V_c_10 nt_c_10 0 0
* Transfer network from port 1 to port 10
R10_1 nt_n_1 nt_c_10 0.003124999999999963
X973 nt_n_1 nt_c_10 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X974 nt_p_1 nt_c_10 rl_admittance res=187800143092.54297 ind=8.409869753766284
X975 nt_p_1 nt_c_10 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X976 nt_p_1 nt_c_10 rl_admittance res=63732557064.23586 ind=35.261662271871394
X977 nt_n_1 nt_c_10 rl_admittance res=112799484372.98152 ind=31.919389834390056
X978 nt_n_1 nt_c_10 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 2 to port 10
R10_2 nt_n_2 nt_c_10 0.003124999999999963
X979 nt_n_2 nt_c_10 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X980 nt_p_2 nt_c_10 rl_admittance res=187800143092.54297 ind=8.409869753766284
X981 nt_p_2 nt_c_10 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X982 nt_p_2 nt_c_10 rl_admittance res=63732557064.23586 ind=35.261662271871394
X983 nt_n_2 nt_c_10 rl_admittance res=112799484372.98152 ind=31.919389834390056
X984 nt_n_2 nt_c_10 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 3 to port 10
R10_3 nt_n_3 nt_c_10 0.003124999999999963
X985 nt_n_3 nt_c_10 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X986 nt_p_3 nt_c_10 rl_admittance res=187800143092.54297 ind=8.409869753766284
X987 nt_p_3 nt_c_10 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X988 nt_p_3 nt_c_10 rl_admittance res=63732557064.23586 ind=35.261662271871394
X989 nt_n_3 nt_c_10 rl_admittance res=112799484372.98152 ind=31.919389834390056
X990 nt_n_3 nt_c_10 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 4 to port 10
R10_4 nt_n_4 nt_c_10 0.003124999999999963
X991 nt_n_4 nt_c_10 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X992 nt_p_4 nt_c_10 rl_admittance res=187800143092.54297 ind=8.409869753766284
X993 nt_p_4 nt_c_10 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X994 nt_p_4 nt_c_10 rl_admittance res=63732557064.23586 ind=35.261662271871394
X995 nt_n_4 nt_c_10 rl_admittance res=112799484372.98152 ind=31.919389834390056
X996 nt_n_4 nt_c_10 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 5 to port 10
R10_5 nt_n_5 nt_c_10 0.003124999999999963
X997 nt_n_5 nt_c_10 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X998 nt_p_5 nt_c_10 rl_admittance res=187800143092.54297 ind=8.409869753766284
X999 nt_p_5 nt_c_10 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1000 nt_p_5 nt_c_10 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1001 nt_n_5 nt_c_10 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1002 nt_n_5 nt_c_10 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 6 to port 10
R10_6 nt_n_6 nt_c_10 0.003124999999999963
X1003 nt_n_6 nt_c_10 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1004 nt_p_6 nt_c_10 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1005 nt_p_6 nt_c_10 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1006 nt_p_6 nt_c_10 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1007 nt_n_6 nt_c_10 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1008 nt_n_6 nt_c_10 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 7 to port 10
R10_7 nt_n_7 nt_c_10 0.003124999999999963
X1009 nt_n_7 nt_c_10 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1010 nt_p_7 nt_c_10 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1011 nt_p_7 nt_c_10 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1012 nt_p_7 nt_c_10 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1013 nt_n_7 nt_c_10 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1014 nt_n_7 nt_c_10 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 8 to port 10
R10_8 nt_n_8 nt_c_10 0.003124999999999963
X1015 nt_n_8 nt_c_10 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1016 nt_p_8 nt_c_10 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1017 nt_p_8 nt_c_10 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1018 nt_p_8 nt_c_10 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1019 nt_n_8 nt_c_10 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1020 nt_n_8 nt_c_10 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 9 to port 10
R10_9 nt_n_9 nt_c_10 0.003124999999999963
X1021 nt_n_9 nt_c_10 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1022 nt_p_9 nt_c_10 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1023 nt_p_9 nt_c_10 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1024 nt_p_9 nt_c_10 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1025 nt_n_9 nt_c_10 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1026 nt_n_9 nt_c_10 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 10 to port 10
R10_10 nt_p_10 nt_c_10 0.0007564900050830436
X1027 nt_p_10 nt_c_10 rl_admittance res=6.713812060922877e+16 ind=0.01239433452121846
X1028 nt_n_10 nt_c_10 rl_admittance res=0.00045787217518182793 ind=2.0503953265122565e-14
X1029 nt_p_10 nt_c_10 rl_admittance res=0.00054254751817662 ind=7.679384261163742e-14
X1030 nt_p_10 nt_c_10 rl_admittance res=0.0005564228350387422 ind=3.0785512135842906e-13
X1031 nt_n_10 nt_c_10 rl_admittance res=0.0005055304090704312 ind=1.4305226916553906e-13
X1032 nt_n_10 nt_c_10 rl_admittance res=0.00047272890640632993 ind=8.643258284073119e-13
* Transfer network from port 11 to port 10
R10_11 nt_n_11 nt_c_10 0.003124999999999963
X1033 nt_n_11 nt_c_10 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1034 nt_p_11 nt_c_10 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1035 nt_p_11 nt_c_10 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1036 nt_p_11 nt_c_10 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1037 nt_n_11 nt_c_10 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1038 nt_n_11 nt_c_10 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 12 to port 10
R10_12 nt_n_12 nt_c_10 0.003124999999999963
X1039 nt_n_12 nt_c_10 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1040 nt_p_12 nt_c_10 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1041 nt_p_12 nt_c_10 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1042 nt_p_12 nt_c_10 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1043 nt_n_12 nt_c_10 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1044 nt_n_12 nt_c_10 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 13 to port 10
R10_13 nt_n_13 nt_c_10 0.003124999999999963
X1045 nt_n_13 nt_c_10 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1046 nt_p_13 nt_c_10 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1047 nt_p_13 nt_c_10 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1048 nt_p_13 nt_c_10 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1049 nt_n_13 nt_c_10 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1050 nt_n_13 nt_c_10 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 14 to port 10
R10_14 nt_n_14 nt_c_10 0.003124999999999963
X1051 nt_n_14 nt_c_10 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1052 nt_p_14 nt_c_10 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1053 nt_p_14 nt_c_10 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1054 nt_p_14 nt_c_10 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1055 nt_n_14 nt_c_10 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1056 nt_n_14 nt_c_10 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 15 to port 10
R10_15 nt_n_15 nt_c_10 0.003124999999999963
X1057 nt_n_15 nt_c_10 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1058 nt_p_15 nt_c_10 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1059 nt_p_15 nt_c_10 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1060 nt_p_15 nt_c_10 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1061 nt_n_15 nt_c_10 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1062 nt_n_15 nt_c_10 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 16 to port 10
R10_16 nt_n_16 nt_c_10 0.003124999999999963
X1063 nt_n_16 nt_c_10 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1064 nt_p_16 nt_c_10 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1065 nt_p_16 nt_c_10 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1066 nt_p_16 nt_c_10 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1067 nt_n_16 nt_c_10 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1068 nt_n_16 nt_c_10 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 17 to port 10
R10_17 nt_n_17 nt_c_10 0.003124999999999963
X1069 nt_n_17 nt_c_10 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1070 nt_p_17 nt_c_10 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1071 nt_p_17 nt_c_10 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1072 nt_p_17 nt_c_10 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1073 nt_n_17 nt_c_10 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1074 nt_n_17 nt_c_10 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 18 to port 10
R10_18 nt_n_18 nt_c_10 0.003124999999999963
X1075 nt_n_18 nt_c_10 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1076 nt_p_18 nt_c_10 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1077 nt_p_18 nt_c_10 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1078 nt_p_18 nt_c_10 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1079 nt_n_18 nt_c_10 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1080 nt_n_18 nt_c_10 rl_admittance res=51262611157.92125 ind=93.72728905498322

* Port network for port 11
R_ref_11 p11 a11 50.0
H_b_11 a11 0 V_c_11 14.142135623730951
* Differential incident wave a sources for transfer from port 11
H_p_11 nt_p_11 nts_p_11 H_b_11 3.5355339059327378
E_p_11 nts_p_11 0 p11 0 0.07071067811865475
E_n_11 0 nt_n_11 nt_p_11 0 1
* Current sensor on center node for transfer to port 11
V_c_11 nt_c_11 0 0
* Transfer network from port 1 to port 11
R11_1 nt_n_1 nt_c_11 0.003124999999999963
X1081 nt_n_1 nt_c_11 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1082 nt_p_1 nt_c_11 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1083 nt_p_1 nt_c_11 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1084 nt_p_1 nt_c_11 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1085 nt_n_1 nt_c_11 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1086 nt_n_1 nt_c_11 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 2 to port 11
R11_2 nt_n_2 nt_c_11 0.003124999999999963
X1087 nt_n_2 nt_c_11 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1088 nt_p_2 nt_c_11 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1089 nt_p_2 nt_c_11 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1090 nt_p_2 nt_c_11 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1091 nt_n_2 nt_c_11 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1092 nt_n_2 nt_c_11 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 3 to port 11
R11_3 nt_n_3 nt_c_11 0.003124999999999963
X1093 nt_n_3 nt_c_11 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1094 nt_p_3 nt_c_11 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1095 nt_p_3 nt_c_11 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1096 nt_p_3 nt_c_11 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1097 nt_n_3 nt_c_11 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1098 nt_n_3 nt_c_11 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 4 to port 11
R11_4 nt_n_4 nt_c_11 0.003124999999999963
X1099 nt_n_4 nt_c_11 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1100 nt_p_4 nt_c_11 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1101 nt_p_4 nt_c_11 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1102 nt_p_4 nt_c_11 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1103 nt_n_4 nt_c_11 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1104 nt_n_4 nt_c_11 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 5 to port 11
R11_5 nt_n_5 nt_c_11 0.003124999999999963
X1105 nt_n_5 nt_c_11 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1106 nt_p_5 nt_c_11 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1107 nt_p_5 nt_c_11 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1108 nt_p_5 nt_c_11 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1109 nt_n_5 nt_c_11 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1110 nt_n_5 nt_c_11 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 6 to port 11
R11_6 nt_n_6 nt_c_11 0.003124999999999963
X1111 nt_n_6 nt_c_11 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1112 nt_p_6 nt_c_11 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1113 nt_p_6 nt_c_11 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1114 nt_p_6 nt_c_11 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1115 nt_n_6 nt_c_11 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1116 nt_n_6 nt_c_11 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 7 to port 11
R11_7 nt_n_7 nt_c_11 0.003124999999999963
X1117 nt_n_7 nt_c_11 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1118 nt_p_7 nt_c_11 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1119 nt_p_7 nt_c_11 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1120 nt_p_7 nt_c_11 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1121 nt_n_7 nt_c_11 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1122 nt_n_7 nt_c_11 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 8 to port 11
R11_8 nt_n_8 nt_c_11 0.003124999999999963
X1123 nt_n_8 nt_c_11 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1124 nt_p_8 nt_c_11 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1125 nt_p_8 nt_c_11 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1126 nt_p_8 nt_c_11 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1127 nt_n_8 nt_c_11 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1128 nt_n_8 nt_c_11 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 9 to port 11
R11_9 nt_n_9 nt_c_11 0.003124999999999963
X1129 nt_n_9 nt_c_11 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1130 nt_p_9 nt_c_11 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1131 nt_p_9 nt_c_11 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1132 nt_p_9 nt_c_11 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1133 nt_n_9 nt_c_11 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1134 nt_n_9 nt_c_11 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 10 to port 11
R11_10 nt_n_10 nt_c_11 0.003124999999999963
X1135 nt_n_10 nt_c_11 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1136 nt_p_10 nt_c_11 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1137 nt_p_10 nt_c_11 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1138 nt_p_10 nt_c_11 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1139 nt_n_10 nt_c_11 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1140 nt_n_10 nt_c_11 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 11 to port 11
R11_11 nt_p_11 nt_c_11 0.0007564900050830436
X1141 nt_p_11 nt_c_11 rl_admittance res=6.713812060922877e+16 ind=0.01239433452121846
X1142 nt_n_11 nt_c_11 rl_admittance res=0.00045787217518182793 ind=2.0503953265122565e-14
X1143 nt_p_11 nt_c_11 rl_admittance res=0.00054254751817662 ind=7.679384261163742e-14
X1144 nt_p_11 nt_c_11 rl_admittance res=0.0005564228350387422 ind=3.0785512135842906e-13
X1145 nt_n_11 nt_c_11 rl_admittance res=0.0005055304090704312 ind=1.4305226916553906e-13
X1146 nt_n_11 nt_c_11 rl_admittance res=0.00047272890640632993 ind=8.643258284073119e-13
* Transfer network from port 12 to port 11
R11_12 nt_n_12 nt_c_11 0.003124999999999963
X1147 nt_n_12 nt_c_11 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1148 nt_p_12 nt_c_11 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1149 nt_p_12 nt_c_11 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1150 nt_p_12 nt_c_11 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1151 nt_n_12 nt_c_11 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1152 nt_n_12 nt_c_11 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 13 to port 11
R11_13 nt_n_13 nt_c_11 0.003124999999999963
X1153 nt_n_13 nt_c_11 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1154 nt_p_13 nt_c_11 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1155 nt_p_13 nt_c_11 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1156 nt_p_13 nt_c_11 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1157 nt_n_13 nt_c_11 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1158 nt_n_13 nt_c_11 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 14 to port 11
R11_14 nt_n_14 nt_c_11 0.003124999999999963
X1159 nt_n_14 nt_c_11 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1160 nt_p_14 nt_c_11 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1161 nt_p_14 nt_c_11 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1162 nt_p_14 nt_c_11 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1163 nt_n_14 nt_c_11 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1164 nt_n_14 nt_c_11 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 15 to port 11
R11_15 nt_n_15 nt_c_11 0.003124999999999963
X1165 nt_n_15 nt_c_11 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1166 nt_p_15 nt_c_11 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1167 nt_p_15 nt_c_11 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1168 nt_p_15 nt_c_11 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1169 nt_n_15 nt_c_11 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1170 nt_n_15 nt_c_11 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 16 to port 11
R11_16 nt_n_16 nt_c_11 0.003124999999999963
X1171 nt_n_16 nt_c_11 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1172 nt_p_16 nt_c_11 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1173 nt_p_16 nt_c_11 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1174 nt_p_16 nt_c_11 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1175 nt_n_16 nt_c_11 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1176 nt_n_16 nt_c_11 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 17 to port 11
R11_17 nt_n_17 nt_c_11 0.003124999999999963
X1177 nt_n_17 nt_c_11 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1178 nt_p_17 nt_c_11 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1179 nt_p_17 nt_c_11 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1180 nt_p_17 nt_c_11 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1181 nt_n_17 nt_c_11 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1182 nt_n_17 nt_c_11 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 18 to port 11
R11_18 nt_n_18 nt_c_11 0.003124999999999963
X1183 nt_n_18 nt_c_11 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1184 nt_p_18 nt_c_11 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1185 nt_p_18 nt_c_11 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1186 nt_p_18 nt_c_11 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1187 nt_n_18 nt_c_11 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1188 nt_n_18 nt_c_11 rl_admittance res=51262611157.92125 ind=93.72728905498322

* Port network for port 12
R_ref_12 p12 a12 50.0
H_b_12 a12 0 V_c_12 14.142135623730951
* Differential incident wave a sources for transfer from port 12
H_p_12 nt_p_12 nts_p_12 H_b_12 3.5355339059327378
E_p_12 nts_p_12 0 p12 0 0.07071067811865475
E_n_12 0 nt_n_12 nt_p_12 0 1
* Current sensor on center node for transfer to port 12
V_c_12 nt_c_12 0 0
* Transfer network from port 1 to port 12
R12_1 nt_n_1 nt_c_12 0.003124999999999963
X1189 nt_n_1 nt_c_12 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1190 nt_p_1 nt_c_12 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1191 nt_p_1 nt_c_12 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1192 nt_p_1 nt_c_12 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1193 nt_n_1 nt_c_12 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1194 nt_n_1 nt_c_12 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 2 to port 12
R12_2 nt_n_2 nt_c_12 0.003124999999999963
X1195 nt_n_2 nt_c_12 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1196 nt_p_2 nt_c_12 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1197 nt_p_2 nt_c_12 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1198 nt_p_2 nt_c_12 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1199 nt_n_2 nt_c_12 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1200 nt_n_2 nt_c_12 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 3 to port 12
R12_3 nt_n_3 nt_c_12 0.003124999999999963
X1201 nt_n_3 nt_c_12 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1202 nt_p_3 nt_c_12 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1203 nt_p_3 nt_c_12 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1204 nt_p_3 nt_c_12 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1205 nt_n_3 nt_c_12 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1206 nt_n_3 nt_c_12 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 4 to port 12
R12_4 nt_n_4 nt_c_12 0.003124999999999963
X1207 nt_n_4 nt_c_12 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1208 nt_p_4 nt_c_12 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1209 nt_p_4 nt_c_12 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1210 nt_p_4 nt_c_12 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1211 nt_n_4 nt_c_12 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1212 nt_n_4 nt_c_12 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 5 to port 12
R12_5 nt_n_5 nt_c_12 0.003124999999999963
X1213 nt_n_5 nt_c_12 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1214 nt_p_5 nt_c_12 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1215 nt_p_5 nt_c_12 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1216 nt_p_5 nt_c_12 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1217 nt_n_5 nt_c_12 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1218 nt_n_5 nt_c_12 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 6 to port 12
R12_6 nt_n_6 nt_c_12 0.003124999999999963
X1219 nt_n_6 nt_c_12 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1220 nt_p_6 nt_c_12 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1221 nt_p_6 nt_c_12 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1222 nt_p_6 nt_c_12 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1223 nt_n_6 nt_c_12 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1224 nt_n_6 nt_c_12 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 7 to port 12
R12_7 nt_n_7 nt_c_12 0.003124999999999963
X1225 nt_n_7 nt_c_12 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1226 nt_p_7 nt_c_12 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1227 nt_p_7 nt_c_12 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1228 nt_p_7 nt_c_12 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1229 nt_n_7 nt_c_12 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1230 nt_n_7 nt_c_12 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 8 to port 12
R12_8 nt_n_8 nt_c_12 0.003124999999999963
X1231 nt_n_8 nt_c_12 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1232 nt_p_8 nt_c_12 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1233 nt_p_8 nt_c_12 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1234 nt_p_8 nt_c_12 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1235 nt_n_8 nt_c_12 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1236 nt_n_8 nt_c_12 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 9 to port 12
R12_9 nt_n_9 nt_c_12 0.003124999999999963
X1237 nt_n_9 nt_c_12 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1238 nt_p_9 nt_c_12 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1239 nt_p_9 nt_c_12 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1240 nt_p_9 nt_c_12 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1241 nt_n_9 nt_c_12 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1242 nt_n_9 nt_c_12 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 10 to port 12
R12_10 nt_n_10 nt_c_12 0.003124999999999963
X1243 nt_n_10 nt_c_12 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1244 nt_p_10 nt_c_12 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1245 nt_p_10 nt_c_12 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1246 nt_p_10 nt_c_12 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1247 nt_n_10 nt_c_12 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1248 nt_n_10 nt_c_12 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 11 to port 12
R12_11 nt_n_11 nt_c_12 0.003124999999999963
X1249 nt_n_11 nt_c_12 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1250 nt_p_11 nt_c_12 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1251 nt_p_11 nt_c_12 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1252 nt_p_11 nt_c_12 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1253 nt_n_11 nt_c_12 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1254 nt_n_11 nt_c_12 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 12 to port 12
R12_12 nt_p_12 nt_c_12 0.0007564900050830436
X1255 nt_p_12 nt_c_12 rl_admittance res=6.713812060922877e+16 ind=0.01239433452121846
X1256 nt_n_12 nt_c_12 rl_admittance res=0.00045787217518182793 ind=2.0503953265122565e-14
X1257 nt_p_12 nt_c_12 rl_admittance res=0.00054254751817662 ind=7.679384261163742e-14
X1258 nt_p_12 nt_c_12 rl_admittance res=0.0005564228350387422 ind=3.0785512135842906e-13
X1259 nt_n_12 nt_c_12 rl_admittance res=0.0005055304090704312 ind=1.4305226916553906e-13
X1260 nt_n_12 nt_c_12 rl_admittance res=0.00047272890640632993 ind=8.643258284073119e-13
* Transfer network from port 13 to port 12
R12_13 nt_n_13 nt_c_12 0.003124999999999963
X1261 nt_n_13 nt_c_12 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1262 nt_p_13 nt_c_12 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1263 nt_p_13 nt_c_12 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1264 nt_p_13 nt_c_12 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1265 nt_n_13 nt_c_12 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1266 nt_n_13 nt_c_12 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 14 to port 12
R12_14 nt_n_14 nt_c_12 0.003124999999999963
X1267 nt_n_14 nt_c_12 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1268 nt_p_14 nt_c_12 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1269 nt_p_14 nt_c_12 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1270 nt_p_14 nt_c_12 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1271 nt_n_14 nt_c_12 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1272 nt_n_14 nt_c_12 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 15 to port 12
R12_15 nt_n_15 nt_c_12 0.003124999999999963
X1273 nt_n_15 nt_c_12 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1274 nt_p_15 nt_c_12 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1275 nt_p_15 nt_c_12 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1276 nt_p_15 nt_c_12 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1277 nt_n_15 nt_c_12 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1278 nt_n_15 nt_c_12 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 16 to port 12
R12_16 nt_n_16 nt_c_12 0.003124999999999963
X1279 nt_n_16 nt_c_12 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1280 nt_p_16 nt_c_12 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1281 nt_p_16 nt_c_12 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1282 nt_p_16 nt_c_12 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1283 nt_n_16 nt_c_12 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1284 nt_n_16 nt_c_12 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 17 to port 12
R12_17 nt_n_17 nt_c_12 0.003124999999999963
X1285 nt_n_17 nt_c_12 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1286 nt_p_17 nt_c_12 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1287 nt_p_17 nt_c_12 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1288 nt_p_17 nt_c_12 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1289 nt_n_17 nt_c_12 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1290 nt_n_17 nt_c_12 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 18 to port 12
R12_18 nt_n_18 nt_c_12 0.003124999999999963
X1291 nt_n_18 nt_c_12 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1292 nt_p_18 nt_c_12 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1293 nt_p_18 nt_c_12 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1294 nt_p_18 nt_c_12 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1295 nt_n_18 nt_c_12 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1296 nt_n_18 nt_c_12 rl_admittance res=51262611157.92125 ind=93.72728905498322

* Port network for port 13
R_ref_13 p13 a13 50.0
H_b_13 a13 0 V_c_13 14.142135623730951
* Differential incident wave a sources for transfer from port 13
H_p_13 nt_p_13 nts_p_13 H_b_13 3.5355339059327378
E_p_13 nts_p_13 0 p13 0 0.07071067811865475
E_n_13 0 nt_n_13 nt_p_13 0 1
* Current sensor on center node for transfer to port 13
V_c_13 nt_c_13 0 0
* Transfer network from port 1 to port 13
R13_1 nt_n_1 nt_c_13 0.003124999999999963
X1297 nt_n_1 nt_c_13 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1298 nt_p_1 nt_c_13 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1299 nt_p_1 nt_c_13 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1300 nt_p_1 nt_c_13 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1301 nt_n_1 nt_c_13 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1302 nt_n_1 nt_c_13 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 2 to port 13
R13_2 nt_n_2 nt_c_13 0.003124999999999963
X1303 nt_n_2 nt_c_13 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1304 nt_p_2 nt_c_13 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1305 nt_p_2 nt_c_13 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1306 nt_p_2 nt_c_13 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1307 nt_n_2 nt_c_13 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1308 nt_n_2 nt_c_13 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 3 to port 13
R13_3 nt_n_3 nt_c_13 0.003124999999999963
X1309 nt_n_3 nt_c_13 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1310 nt_p_3 nt_c_13 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1311 nt_p_3 nt_c_13 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1312 nt_p_3 nt_c_13 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1313 nt_n_3 nt_c_13 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1314 nt_n_3 nt_c_13 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 4 to port 13
R13_4 nt_n_4 nt_c_13 0.003124999999999963
X1315 nt_n_4 nt_c_13 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1316 nt_p_4 nt_c_13 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1317 nt_p_4 nt_c_13 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1318 nt_p_4 nt_c_13 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1319 nt_n_4 nt_c_13 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1320 nt_n_4 nt_c_13 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 5 to port 13
R13_5 nt_n_5 nt_c_13 0.003124999999999963
X1321 nt_n_5 nt_c_13 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1322 nt_p_5 nt_c_13 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1323 nt_p_5 nt_c_13 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1324 nt_p_5 nt_c_13 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1325 nt_n_5 nt_c_13 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1326 nt_n_5 nt_c_13 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 6 to port 13
R13_6 nt_n_6 nt_c_13 0.003124999999999963
X1327 nt_n_6 nt_c_13 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1328 nt_p_6 nt_c_13 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1329 nt_p_6 nt_c_13 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1330 nt_p_6 nt_c_13 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1331 nt_n_6 nt_c_13 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1332 nt_n_6 nt_c_13 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 7 to port 13
R13_7 nt_n_7 nt_c_13 0.003124999999999963
X1333 nt_n_7 nt_c_13 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1334 nt_p_7 nt_c_13 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1335 nt_p_7 nt_c_13 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1336 nt_p_7 nt_c_13 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1337 nt_n_7 nt_c_13 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1338 nt_n_7 nt_c_13 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 8 to port 13
R13_8 nt_n_8 nt_c_13 0.003124999999999963
X1339 nt_n_8 nt_c_13 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1340 nt_p_8 nt_c_13 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1341 nt_p_8 nt_c_13 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1342 nt_p_8 nt_c_13 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1343 nt_n_8 nt_c_13 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1344 nt_n_8 nt_c_13 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 9 to port 13
R13_9 nt_n_9 nt_c_13 0.003124999999999963
X1345 nt_n_9 nt_c_13 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1346 nt_p_9 nt_c_13 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1347 nt_p_9 nt_c_13 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1348 nt_p_9 nt_c_13 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1349 nt_n_9 nt_c_13 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1350 nt_n_9 nt_c_13 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 10 to port 13
R13_10 nt_n_10 nt_c_13 0.003124999999999963
X1351 nt_n_10 nt_c_13 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1352 nt_p_10 nt_c_13 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1353 nt_p_10 nt_c_13 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1354 nt_p_10 nt_c_13 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1355 nt_n_10 nt_c_13 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1356 nt_n_10 nt_c_13 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 11 to port 13
R13_11 nt_n_11 nt_c_13 0.003124999999999963
X1357 nt_n_11 nt_c_13 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1358 nt_p_11 nt_c_13 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1359 nt_p_11 nt_c_13 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1360 nt_p_11 nt_c_13 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1361 nt_n_11 nt_c_13 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1362 nt_n_11 nt_c_13 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 12 to port 13
R13_12 nt_n_12 nt_c_13 0.003124999999999963
X1363 nt_n_12 nt_c_13 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1364 nt_p_12 nt_c_13 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1365 nt_p_12 nt_c_13 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1366 nt_p_12 nt_c_13 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1367 nt_n_12 nt_c_13 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1368 nt_n_12 nt_c_13 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 13 to port 13
R13_13 nt_p_13 nt_c_13 0.0007564900050830436
X1369 nt_p_13 nt_c_13 rl_admittance res=6.713812060922877e+16 ind=0.01239433452121846
X1370 nt_n_13 nt_c_13 rl_admittance res=0.00045787217518182793 ind=2.0503953265122565e-14
X1371 nt_p_13 nt_c_13 rl_admittance res=0.00054254751817662 ind=7.679384261163742e-14
X1372 nt_p_13 nt_c_13 rl_admittance res=0.0005564228350387422 ind=3.0785512135842906e-13
X1373 nt_n_13 nt_c_13 rl_admittance res=0.0005055304090704312 ind=1.4305226916553906e-13
X1374 nt_n_13 nt_c_13 rl_admittance res=0.00047272890640632993 ind=8.643258284073119e-13
* Transfer network from port 14 to port 13
R13_14 nt_n_14 nt_c_13 0.003124999999999963
X1375 nt_n_14 nt_c_13 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1376 nt_p_14 nt_c_13 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1377 nt_p_14 nt_c_13 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1378 nt_p_14 nt_c_13 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1379 nt_n_14 nt_c_13 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1380 nt_n_14 nt_c_13 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 15 to port 13
R13_15 nt_n_15 nt_c_13 0.003124999999999963
X1381 nt_n_15 nt_c_13 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1382 nt_p_15 nt_c_13 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1383 nt_p_15 nt_c_13 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1384 nt_p_15 nt_c_13 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1385 nt_n_15 nt_c_13 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1386 nt_n_15 nt_c_13 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 16 to port 13
R13_16 nt_n_16 nt_c_13 0.003124999999999963
X1387 nt_n_16 nt_c_13 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1388 nt_p_16 nt_c_13 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1389 nt_p_16 nt_c_13 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1390 nt_p_16 nt_c_13 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1391 nt_n_16 nt_c_13 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1392 nt_n_16 nt_c_13 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 17 to port 13
R13_17 nt_n_17 nt_c_13 0.003124999999999963
X1393 nt_n_17 nt_c_13 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1394 nt_p_17 nt_c_13 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1395 nt_p_17 nt_c_13 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1396 nt_p_17 nt_c_13 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1397 nt_n_17 nt_c_13 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1398 nt_n_17 nt_c_13 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 18 to port 13
R13_18 nt_n_18 nt_c_13 0.003124999999999963
X1399 nt_n_18 nt_c_13 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1400 nt_p_18 nt_c_13 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1401 nt_p_18 nt_c_13 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1402 nt_p_18 nt_c_13 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1403 nt_n_18 nt_c_13 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1404 nt_n_18 nt_c_13 rl_admittance res=51262611157.92125 ind=93.72728905498322

* Port network for port 14
R_ref_14 p14 a14 50.0
H_b_14 a14 0 V_c_14 14.142135623730951
* Differential incident wave a sources for transfer from port 14
H_p_14 nt_p_14 nts_p_14 H_b_14 3.5355339059327378
E_p_14 nts_p_14 0 p14 0 0.07071067811865475
E_n_14 0 nt_n_14 nt_p_14 0 1
* Current sensor on center node for transfer to port 14
V_c_14 nt_c_14 0 0
* Transfer network from port 1 to port 14
R14_1 nt_n_1 nt_c_14 0.003124999999999963
X1405 nt_n_1 nt_c_14 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1406 nt_p_1 nt_c_14 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1407 nt_p_1 nt_c_14 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1408 nt_p_1 nt_c_14 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1409 nt_n_1 nt_c_14 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1410 nt_n_1 nt_c_14 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 2 to port 14
R14_2 nt_n_2 nt_c_14 0.003124999999999963
X1411 nt_n_2 nt_c_14 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1412 nt_p_2 nt_c_14 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1413 nt_p_2 nt_c_14 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1414 nt_p_2 nt_c_14 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1415 nt_n_2 nt_c_14 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1416 nt_n_2 nt_c_14 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 3 to port 14
R14_3 nt_n_3 nt_c_14 0.003124999999999963
X1417 nt_n_3 nt_c_14 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1418 nt_p_3 nt_c_14 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1419 nt_p_3 nt_c_14 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1420 nt_p_3 nt_c_14 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1421 nt_n_3 nt_c_14 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1422 nt_n_3 nt_c_14 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 4 to port 14
R14_4 nt_n_4 nt_c_14 0.003124999999999963
X1423 nt_n_4 nt_c_14 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1424 nt_p_4 nt_c_14 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1425 nt_p_4 nt_c_14 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1426 nt_p_4 nt_c_14 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1427 nt_n_4 nt_c_14 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1428 nt_n_4 nt_c_14 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 5 to port 14
R14_5 nt_n_5 nt_c_14 0.003124999999999963
X1429 nt_n_5 nt_c_14 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1430 nt_p_5 nt_c_14 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1431 nt_p_5 nt_c_14 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1432 nt_p_5 nt_c_14 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1433 nt_n_5 nt_c_14 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1434 nt_n_5 nt_c_14 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 6 to port 14
R14_6 nt_n_6 nt_c_14 0.003124999999999963
X1435 nt_n_6 nt_c_14 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1436 nt_p_6 nt_c_14 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1437 nt_p_6 nt_c_14 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1438 nt_p_6 nt_c_14 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1439 nt_n_6 nt_c_14 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1440 nt_n_6 nt_c_14 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 7 to port 14
R14_7 nt_n_7 nt_c_14 0.003124999999999963
X1441 nt_n_7 nt_c_14 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1442 nt_p_7 nt_c_14 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1443 nt_p_7 nt_c_14 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1444 nt_p_7 nt_c_14 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1445 nt_n_7 nt_c_14 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1446 nt_n_7 nt_c_14 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 8 to port 14
R14_8 nt_n_8 nt_c_14 0.003124999999999963
X1447 nt_n_8 nt_c_14 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1448 nt_p_8 nt_c_14 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1449 nt_p_8 nt_c_14 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1450 nt_p_8 nt_c_14 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1451 nt_n_8 nt_c_14 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1452 nt_n_8 nt_c_14 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 9 to port 14
R14_9 nt_n_9 nt_c_14 0.003124999999999963
X1453 nt_n_9 nt_c_14 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1454 nt_p_9 nt_c_14 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1455 nt_p_9 nt_c_14 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1456 nt_p_9 nt_c_14 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1457 nt_n_9 nt_c_14 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1458 nt_n_9 nt_c_14 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 10 to port 14
R14_10 nt_n_10 nt_c_14 0.003124999999999963
X1459 nt_n_10 nt_c_14 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1460 nt_p_10 nt_c_14 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1461 nt_p_10 nt_c_14 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1462 nt_p_10 nt_c_14 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1463 nt_n_10 nt_c_14 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1464 nt_n_10 nt_c_14 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 11 to port 14
R14_11 nt_n_11 nt_c_14 0.003124999999999963
X1465 nt_n_11 nt_c_14 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1466 nt_p_11 nt_c_14 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1467 nt_p_11 nt_c_14 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1468 nt_p_11 nt_c_14 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1469 nt_n_11 nt_c_14 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1470 nt_n_11 nt_c_14 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 12 to port 14
R14_12 nt_n_12 nt_c_14 0.003124999999999963
X1471 nt_n_12 nt_c_14 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1472 nt_p_12 nt_c_14 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1473 nt_p_12 nt_c_14 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1474 nt_p_12 nt_c_14 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1475 nt_n_12 nt_c_14 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1476 nt_n_12 nt_c_14 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 13 to port 14
R14_13 nt_n_13 nt_c_14 0.003124999999999963
X1477 nt_n_13 nt_c_14 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1478 nt_p_13 nt_c_14 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1479 nt_p_13 nt_c_14 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1480 nt_p_13 nt_c_14 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1481 nt_n_13 nt_c_14 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1482 nt_n_13 nt_c_14 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 14 to port 14
R14_14 nt_p_14 nt_c_14 0.0007564900050830436
X1483 nt_p_14 nt_c_14 rl_admittance res=6.713812060922877e+16 ind=0.01239433452121846
X1484 nt_n_14 nt_c_14 rl_admittance res=0.00045787217518182793 ind=2.0503953265122565e-14
X1485 nt_p_14 nt_c_14 rl_admittance res=0.00054254751817662 ind=7.679384261163742e-14
X1486 nt_p_14 nt_c_14 rl_admittance res=0.0005564228350387422 ind=3.0785512135842906e-13
X1487 nt_n_14 nt_c_14 rl_admittance res=0.0005055304090704312 ind=1.4305226916553906e-13
X1488 nt_n_14 nt_c_14 rl_admittance res=0.00047272890640632993 ind=8.643258284073119e-13
* Transfer network from port 15 to port 14
R14_15 nt_n_15 nt_c_14 0.003124999999999963
X1489 nt_n_15 nt_c_14 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1490 nt_p_15 nt_c_14 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1491 nt_p_15 nt_c_14 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1492 nt_p_15 nt_c_14 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1493 nt_n_15 nt_c_14 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1494 nt_n_15 nt_c_14 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 16 to port 14
R14_16 nt_n_16 nt_c_14 0.003124999999999963
X1495 nt_n_16 nt_c_14 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1496 nt_p_16 nt_c_14 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1497 nt_p_16 nt_c_14 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1498 nt_p_16 nt_c_14 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1499 nt_n_16 nt_c_14 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1500 nt_n_16 nt_c_14 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 17 to port 14
R14_17 nt_n_17 nt_c_14 0.003124999999999963
X1501 nt_n_17 nt_c_14 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1502 nt_p_17 nt_c_14 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1503 nt_p_17 nt_c_14 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1504 nt_p_17 nt_c_14 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1505 nt_n_17 nt_c_14 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1506 nt_n_17 nt_c_14 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 18 to port 14
R14_18 nt_n_18 nt_c_14 0.003124999999999963
X1507 nt_n_18 nt_c_14 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1508 nt_p_18 nt_c_14 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1509 nt_p_18 nt_c_14 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1510 nt_p_18 nt_c_14 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1511 nt_n_18 nt_c_14 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1512 nt_n_18 nt_c_14 rl_admittance res=51262611157.92125 ind=93.72728905498322

* Port network for port 15
R_ref_15 p15 a15 50.0
H_b_15 a15 0 V_c_15 14.142135623730951
* Differential incident wave a sources for transfer from port 15
H_p_15 nt_p_15 nts_p_15 H_b_15 3.5355339059327378
E_p_15 nts_p_15 0 p15 0 0.07071067811865475
E_n_15 0 nt_n_15 nt_p_15 0 1
* Current sensor on center node for transfer to port 15
V_c_15 nt_c_15 0 0
* Transfer network from port 1 to port 15
R15_1 nt_n_1 nt_c_15 0.003124999999999963
X1513 nt_n_1 nt_c_15 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1514 nt_p_1 nt_c_15 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1515 nt_p_1 nt_c_15 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1516 nt_p_1 nt_c_15 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1517 nt_n_1 nt_c_15 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1518 nt_n_1 nt_c_15 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 2 to port 15
R15_2 nt_n_2 nt_c_15 0.003124999999999963
X1519 nt_n_2 nt_c_15 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1520 nt_p_2 nt_c_15 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1521 nt_p_2 nt_c_15 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1522 nt_p_2 nt_c_15 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1523 nt_n_2 nt_c_15 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1524 nt_n_2 nt_c_15 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 3 to port 15
R15_3 nt_n_3 nt_c_15 0.003124999999999963
X1525 nt_n_3 nt_c_15 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1526 nt_p_3 nt_c_15 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1527 nt_p_3 nt_c_15 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1528 nt_p_3 nt_c_15 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1529 nt_n_3 nt_c_15 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1530 nt_n_3 nt_c_15 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 4 to port 15
R15_4 nt_n_4 nt_c_15 0.003124999999999963
X1531 nt_n_4 nt_c_15 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1532 nt_p_4 nt_c_15 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1533 nt_p_4 nt_c_15 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1534 nt_p_4 nt_c_15 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1535 nt_n_4 nt_c_15 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1536 nt_n_4 nt_c_15 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 5 to port 15
R15_5 nt_n_5 nt_c_15 0.003124999999999963
X1537 nt_n_5 nt_c_15 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1538 nt_p_5 nt_c_15 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1539 nt_p_5 nt_c_15 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1540 nt_p_5 nt_c_15 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1541 nt_n_5 nt_c_15 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1542 nt_n_5 nt_c_15 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 6 to port 15
R15_6 nt_n_6 nt_c_15 0.003124999999999963
X1543 nt_n_6 nt_c_15 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1544 nt_p_6 nt_c_15 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1545 nt_p_6 nt_c_15 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1546 nt_p_6 nt_c_15 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1547 nt_n_6 nt_c_15 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1548 nt_n_6 nt_c_15 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 7 to port 15
R15_7 nt_n_7 nt_c_15 0.003124999999999963
X1549 nt_n_7 nt_c_15 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1550 nt_p_7 nt_c_15 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1551 nt_p_7 nt_c_15 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1552 nt_p_7 nt_c_15 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1553 nt_n_7 nt_c_15 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1554 nt_n_7 nt_c_15 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 8 to port 15
R15_8 nt_n_8 nt_c_15 0.003124999999999963
X1555 nt_n_8 nt_c_15 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1556 nt_p_8 nt_c_15 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1557 nt_p_8 nt_c_15 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1558 nt_p_8 nt_c_15 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1559 nt_n_8 nt_c_15 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1560 nt_n_8 nt_c_15 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 9 to port 15
R15_9 nt_n_9 nt_c_15 0.003124999999999963
X1561 nt_n_9 nt_c_15 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1562 nt_p_9 nt_c_15 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1563 nt_p_9 nt_c_15 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1564 nt_p_9 nt_c_15 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1565 nt_n_9 nt_c_15 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1566 nt_n_9 nt_c_15 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 10 to port 15
R15_10 nt_n_10 nt_c_15 0.003124999999999963
X1567 nt_n_10 nt_c_15 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1568 nt_p_10 nt_c_15 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1569 nt_p_10 nt_c_15 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1570 nt_p_10 nt_c_15 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1571 nt_n_10 nt_c_15 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1572 nt_n_10 nt_c_15 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 11 to port 15
R15_11 nt_n_11 nt_c_15 0.003124999999999963
X1573 nt_n_11 nt_c_15 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1574 nt_p_11 nt_c_15 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1575 nt_p_11 nt_c_15 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1576 nt_p_11 nt_c_15 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1577 nt_n_11 nt_c_15 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1578 nt_n_11 nt_c_15 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 12 to port 15
R15_12 nt_n_12 nt_c_15 0.003124999999999963
X1579 nt_n_12 nt_c_15 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1580 nt_p_12 nt_c_15 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1581 nt_p_12 nt_c_15 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1582 nt_p_12 nt_c_15 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1583 nt_n_12 nt_c_15 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1584 nt_n_12 nt_c_15 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 13 to port 15
R15_13 nt_n_13 nt_c_15 0.003124999999999963
X1585 nt_n_13 nt_c_15 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1586 nt_p_13 nt_c_15 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1587 nt_p_13 nt_c_15 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1588 nt_p_13 nt_c_15 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1589 nt_n_13 nt_c_15 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1590 nt_n_13 nt_c_15 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 14 to port 15
R15_14 nt_n_14 nt_c_15 0.003124999999999963
X1591 nt_n_14 nt_c_15 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1592 nt_p_14 nt_c_15 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1593 nt_p_14 nt_c_15 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1594 nt_p_14 nt_c_15 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1595 nt_n_14 nt_c_15 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1596 nt_n_14 nt_c_15 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 15 to port 15
R15_15 nt_p_15 nt_c_15 0.0007564900050830436
X1597 nt_p_15 nt_c_15 rl_admittance res=6.713812060922877e+16 ind=0.01239433452121846
X1598 nt_n_15 nt_c_15 rl_admittance res=0.00045787217518182793 ind=2.0503953265122565e-14
X1599 nt_p_15 nt_c_15 rl_admittance res=0.00054254751817662 ind=7.679384261163742e-14
X1600 nt_p_15 nt_c_15 rl_admittance res=0.0005564228350387422 ind=3.0785512135842906e-13
X1601 nt_n_15 nt_c_15 rl_admittance res=0.0005055304090704312 ind=1.4305226916553906e-13
X1602 nt_n_15 nt_c_15 rl_admittance res=0.00047272890640632993 ind=8.643258284073119e-13
* Transfer network from port 16 to port 15
R15_16 nt_n_16 nt_c_15 0.003124999999999963
X1603 nt_n_16 nt_c_15 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1604 nt_p_16 nt_c_15 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1605 nt_p_16 nt_c_15 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1606 nt_p_16 nt_c_15 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1607 nt_n_16 nt_c_15 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1608 nt_n_16 nt_c_15 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 17 to port 15
R15_17 nt_n_17 nt_c_15 0.003124999999999963
X1609 nt_n_17 nt_c_15 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1610 nt_p_17 nt_c_15 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1611 nt_p_17 nt_c_15 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1612 nt_p_17 nt_c_15 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1613 nt_n_17 nt_c_15 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1614 nt_n_17 nt_c_15 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 18 to port 15
R15_18 nt_n_18 nt_c_15 0.003124999999999963
X1615 nt_n_18 nt_c_15 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1616 nt_p_18 nt_c_15 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1617 nt_p_18 nt_c_15 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1618 nt_p_18 nt_c_15 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1619 nt_n_18 nt_c_15 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1620 nt_n_18 nt_c_15 rl_admittance res=51262611157.92125 ind=93.72728905498322

* Port network for port 16
R_ref_16 p16 a16 50.0
H_b_16 a16 0 V_c_16 14.142135623730951
* Differential incident wave a sources for transfer from port 16
H_p_16 nt_p_16 nts_p_16 H_b_16 3.5355339059327378
E_p_16 nts_p_16 0 p16 0 0.07071067811865475
E_n_16 0 nt_n_16 nt_p_16 0 1
* Current sensor on center node for transfer to port 16
V_c_16 nt_c_16 0 0
* Transfer network from port 1 to port 16
R16_1 nt_n_1 nt_c_16 0.003124999999999963
X1621 nt_n_1 nt_c_16 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1622 nt_p_1 nt_c_16 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1623 nt_p_1 nt_c_16 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1624 nt_p_1 nt_c_16 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1625 nt_n_1 nt_c_16 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1626 nt_n_1 nt_c_16 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 2 to port 16
R16_2 nt_n_2 nt_c_16 0.003124999999999963
X1627 nt_n_2 nt_c_16 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1628 nt_p_2 nt_c_16 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1629 nt_p_2 nt_c_16 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1630 nt_p_2 nt_c_16 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1631 nt_n_2 nt_c_16 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1632 nt_n_2 nt_c_16 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 3 to port 16
R16_3 nt_n_3 nt_c_16 0.003124999999999963
X1633 nt_n_3 nt_c_16 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1634 nt_p_3 nt_c_16 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1635 nt_p_3 nt_c_16 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1636 nt_p_3 nt_c_16 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1637 nt_n_3 nt_c_16 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1638 nt_n_3 nt_c_16 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 4 to port 16
R16_4 nt_n_4 nt_c_16 0.003124999999999963
X1639 nt_n_4 nt_c_16 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1640 nt_p_4 nt_c_16 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1641 nt_p_4 nt_c_16 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1642 nt_p_4 nt_c_16 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1643 nt_n_4 nt_c_16 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1644 nt_n_4 nt_c_16 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 5 to port 16
R16_5 nt_n_5 nt_c_16 0.003124999999999963
X1645 nt_n_5 nt_c_16 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1646 nt_p_5 nt_c_16 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1647 nt_p_5 nt_c_16 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1648 nt_p_5 nt_c_16 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1649 nt_n_5 nt_c_16 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1650 nt_n_5 nt_c_16 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 6 to port 16
R16_6 nt_n_6 nt_c_16 0.003124999999999963
X1651 nt_n_6 nt_c_16 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1652 nt_p_6 nt_c_16 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1653 nt_p_6 nt_c_16 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1654 nt_p_6 nt_c_16 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1655 nt_n_6 nt_c_16 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1656 nt_n_6 nt_c_16 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 7 to port 16
R16_7 nt_n_7 nt_c_16 0.003124999999999963
X1657 nt_n_7 nt_c_16 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1658 nt_p_7 nt_c_16 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1659 nt_p_7 nt_c_16 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1660 nt_p_7 nt_c_16 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1661 nt_n_7 nt_c_16 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1662 nt_n_7 nt_c_16 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 8 to port 16
R16_8 nt_n_8 nt_c_16 0.003124999999999963
X1663 nt_n_8 nt_c_16 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1664 nt_p_8 nt_c_16 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1665 nt_p_8 nt_c_16 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1666 nt_p_8 nt_c_16 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1667 nt_n_8 nt_c_16 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1668 nt_n_8 nt_c_16 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 9 to port 16
R16_9 nt_n_9 nt_c_16 0.003124999999999963
X1669 nt_n_9 nt_c_16 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1670 nt_p_9 nt_c_16 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1671 nt_p_9 nt_c_16 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1672 nt_p_9 nt_c_16 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1673 nt_n_9 nt_c_16 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1674 nt_n_9 nt_c_16 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 10 to port 16
R16_10 nt_n_10 nt_c_16 0.003124999999999963
X1675 nt_n_10 nt_c_16 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1676 nt_p_10 nt_c_16 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1677 nt_p_10 nt_c_16 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1678 nt_p_10 nt_c_16 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1679 nt_n_10 nt_c_16 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1680 nt_n_10 nt_c_16 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 11 to port 16
R16_11 nt_n_11 nt_c_16 0.003124999999999963
X1681 nt_n_11 nt_c_16 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1682 nt_p_11 nt_c_16 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1683 nt_p_11 nt_c_16 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1684 nt_p_11 nt_c_16 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1685 nt_n_11 nt_c_16 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1686 nt_n_11 nt_c_16 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 12 to port 16
R16_12 nt_n_12 nt_c_16 0.003124999999999963
X1687 nt_n_12 nt_c_16 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1688 nt_p_12 nt_c_16 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1689 nt_p_12 nt_c_16 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1690 nt_p_12 nt_c_16 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1691 nt_n_12 nt_c_16 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1692 nt_n_12 nt_c_16 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 13 to port 16
R16_13 nt_n_13 nt_c_16 0.003124999999999963
X1693 nt_n_13 nt_c_16 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1694 nt_p_13 nt_c_16 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1695 nt_p_13 nt_c_16 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1696 nt_p_13 nt_c_16 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1697 nt_n_13 nt_c_16 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1698 nt_n_13 nt_c_16 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 14 to port 16
R16_14 nt_n_14 nt_c_16 0.003124999999999963
X1699 nt_n_14 nt_c_16 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1700 nt_p_14 nt_c_16 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1701 nt_p_14 nt_c_16 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1702 nt_p_14 nt_c_16 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1703 nt_n_14 nt_c_16 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1704 nt_n_14 nt_c_16 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 15 to port 16
R16_15 nt_n_15 nt_c_16 0.003124999999999963
X1705 nt_n_15 nt_c_16 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1706 nt_p_15 nt_c_16 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1707 nt_p_15 nt_c_16 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1708 nt_p_15 nt_c_16 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1709 nt_n_15 nt_c_16 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1710 nt_n_15 nt_c_16 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 16 to port 16
R16_16 nt_p_16 nt_c_16 0.0007564900050830436
X1711 nt_p_16 nt_c_16 rl_admittance res=6.713812060922877e+16 ind=0.01239433452121846
X1712 nt_n_16 nt_c_16 rl_admittance res=0.00045787217518182793 ind=2.0503953265122565e-14
X1713 nt_p_16 nt_c_16 rl_admittance res=0.00054254751817662 ind=7.679384261163742e-14
X1714 nt_p_16 nt_c_16 rl_admittance res=0.0005564228350387422 ind=3.0785512135842906e-13
X1715 nt_n_16 nt_c_16 rl_admittance res=0.0005055304090704312 ind=1.4305226916553906e-13
X1716 nt_n_16 nt_c_16 rl_admittance res=0.00047272890640632993 ind=8.643258284073119e-13
* Transfer network from port 17 to port 16
R16_17 nt_n_17 nt_c_16 0.003124999999999963
X1717 nt_n_17 nt_c_16 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1718 nt_p_17 nt_c_16 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1719 nt_p_17 nt_c_16 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1720 nt_p_17 nt_c_16 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1721 nt_n_17 nt_c_16 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1722 nt_n_17 nt_c_16 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 18 to port 16
R16_18 nt_n_18 nt_c_16 0.003124999999999963
X1723 nt_n_18 nt_c_16 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1724 nt_p_18 nt_c_16 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1725 nt_p_18 nt_c_16 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1726 nt_p_18 nt_c_16 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1727 nt_n_18 nt_c_16 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1728 nt_n_18 nt_c_16 rl_admittance res=51262611157.92125 ind=93.72728905498322

* Port network for port 17
R_ref_17 p17 a17 50.0
H_b_17 a17 0 V_c_17 14.142135623730951
* Differential incident wave a sources for transfer from port 17
H_p_17 nt_p_17 nts_p_17 H_b_17 3.5355339059327378
E_p_17 nts_p_17 0 p17 0 0.07071067811865475
E_n_17 0 nt_n_17 nt_p_17 0 1
* Current sensor on center node for transfer to port 17
V_c_17 nt_c_17 0 0
* Transfer network from port 1 to port 17
R17_1 nt_n_1 nt_c_17 0.003124999999999963
X1729 nt_n_1 nt_c_17 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1730 nt_p_1 nt_c_17 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1731 nt_p_1 nt_c_17 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1732 nt_p_1 nt_c_17 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1733 nt_n_1 nt_c_17 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1734 nt_n_1 nt_c_17 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 2 to port 17
R17_2 nt_n_2 nt_c_17 0.003124999999999963
X1735 nt_n_2 nt_c_17 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1736 nt_p_2 nt_c_17 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1737 nt_p_2 nt_c_17 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1738 nt_p_2 nt_c_17 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1739 nt_n_2 nt_c_17 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1740 nt_n_2 nt_c_17 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 3 to port 17
R17_3 nt_n_3 nt_c_17 0.003124999999999963
X1741 nt_n_3 nt_c_17 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1742 nt_p_3 nt_c_17 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1743 nt_p_3 nt_c_17 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1744 nt_p_3 nt_c_17 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1745 nt_n_3 nt_c_17 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1746 nt_n_3 nt_c_17 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 4 to port 17
R17_4 nt_n_4 nt_c_17 0.003124999999999963
X1747 nt_n_4 nt_c_17 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1748 nt_p_4 nt_c_17 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1749 nt_p_4 nt_c_17 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1750 nt_p_4 nt_c_17 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1751 nt_n_4 nt_c_17 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1752 nt_n_4 nt_c_17 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 5 to port 17
R17_5 nt_n_5 nt_c_17 0.003124999999999963
X1753 nt_n_5 nt_c_17 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1754 nt_p_5 nt_c_17 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1755 nt_p_5 nt_c_17 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1756 nt_p_5 nt_c_17 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1757 nt_n_5 nt_c_17 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1758 nt_n_5 nt_c_17 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 6 to port 17
R17_6 nt_n_6 nt_c_17 0.003124999999999963
X1759 nt_n_6 nt_c_17 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1760 nt_p_6 nt_c_17 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1761 nt_p_6 nt_c_17 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1762 nt_p_6 nt_c_17 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1763 nt_n_6 nt_c_17 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1764 nt_n_6 nt_c_17 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 7 to port 17
R17_7 nt_n_7 nt_c_17 0.003124999999999963
X1765 nt_n_7 nt_c_17 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1766 nt_p_7 nt_c_17 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1767 nt_p_7 nt_c_17 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1768 nt_p_7 nt_c_17 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1769 nt_n_7 nt_c_17 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1770 nt_n_7 nt_c_17 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 8 to port 17
R17_8 nt_n_8 nt_c_17 0.003124999999999963
X1771 nt_n_8 nt_c_17 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1772 nt_p_8 nt_c_17 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1773 nt_p_8 nt_c_17 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1774 nt_p_8 nt_c_17 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1775 nt_n_8 nt_c_17 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1776 nt_n_8 nt_c_17 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 9 to port 17
R17_9 nt_n_9 nt_c_17 0.003124999999999963
X1777 nt_n_9 nt_c_17 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1778 nt_p_9 nt_c_17 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1779 nt_p_9 nt_c_17 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1780 nt_p_9 nt_c_17 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1781 nt_n_9 nt_c_17 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1782 nt_n_9 nt_c_17 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 10 to port 17
R17_10 nt_n_10 nt_c_17 0.003124999999999963
X1783 nt_n_10 nt_c_17 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1784 nt_p_10 nt_c_17 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1785 nt_p_10 nt_c_17 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1786 nt_p_10 nt_c_17 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1787 nt_n_10 nt_c_17 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1788 nt_n_10 nt_c_17 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 11 to port 17
R17_11 nt_n_11 nt_c_17 0.003124999999999963
X1789 nt_n_11 nt_c_17 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1790 nt_p_11 nt_c_17 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1791 nt_p_11 nt_c_17 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1792 nt_p_11 nt_c_17 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1793 nt_n_11 nt_c_17 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1794 nt_n_11 nt_c_17 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 12 to port 17
R17_12 nt_n_12 nt_c_17 0.003124999999999963
X1795 nt_n_12 nt_c_17 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1796 nt_p_12 nt_c_17 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1797 nt_p_12 nt_c_17 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1798 nt_p_12 nt_c_17 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1799 nt_n_12 nt_c_17 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1800 nt_n_12 nt_c_17 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 13 to port 17
R17_13 nt_n_13 nt_c_17 0.003124999999999963
X1801 nt_n_13 nt_c_17 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1802 nt_p_13 nt_c_17 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1803 nt_p_13 nt_c_17 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1804 nt_p_13 nt_c_17 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1805 nt_n_13 nt_c_17 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1806 nt_n_13 nt_c_17 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 14 to port 17
R17_14 nt_n_14 nt_c_17 0.003124999999999963
X1807 nt_n_14 nt_c_17 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1808 nt_p_14 nt_c_17 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1809 nt_p_14 nt_c_17 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1810 nt_p_14 nt_c_17 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1811 nt_n_14 nt_c_17 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1812 nt_n_14 nt_c_17 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 15 to port 17
R17_15 nt_n_15 nt_c_17 0.003124999999999963
X1813 nt_n_15 nt_c_17 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1814 nt_p_15 nt_c_17 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1815 nt_p_15 nt_c_17 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1816 nt_p_15 nt_c_17 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1817 nt_n_15 nt_c_17 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1818 nt_n_15 nt_c_17 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 16 to port 17
R17_16 nt_n_16 nt_c_17 0.003124999999999963
X1819 nt_n_16 nt_c_17 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1820 nt_p_16 nt_c_17 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1821 nt_p_16 nt_c_17 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1822 nt_p_16 nt_c_17 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1823 nt_n_16 nt_c_17 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1824 nt_n_16 nt_c_17 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 17 to port 17
R17_17 nt_p_17 nt_c_17 0.0007564900050830436
X1825 nt_p_17 nt_c_17 rl_admittance res=6.713812060922877e+16 ind=0.01239433452121846
X1826 nt_n_17 nt_c_17 rl_admittance res=0.00045787217518182793 ind=2.0503953265122565e-14
X1827 nt_p_17 nt_c_17 rl_admittance res=0.00054254751817662 ind=7.679384261163742e-14
X1828 nt_p_17 nt_c_17 rl_admittance res=0.0005564228350387422 ind=3.0785512135842906e-13
X1829 nt_n_17 nt_c_17 rl_admittance res=0.0005055304090704312 ind=1.4305226916553906e-13
X1830 nt_n_17 nt_c_17 rl_admittance res=0.00047272890640632993 ind=8.643258284073119e-13
* Transfer network from port 18 to port 17
R17_18 nt_n_18 nt_c_17 0.003124999999999963
X1831 nt_n_18 nt_c_17 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1832 nt_p_18 nt_c_17 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1833 nt_p_18 nt_c_17 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1834 nt_p_18 nt_c_17 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1835 nt_n_18 nt_c_17 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1836 nt_n_18 nt_c_17 rl_admittance res=51262611157.92125 ind=93.72728905498322

* Port network for port 18
R_ref_18 p18 a18 50.0
H_b_18 a18 0 V_c_18 14.142135623730951
* Differential incident wave a sources for transfer from port 18
H_p_18 nt_p_18 nts_p_18 H_b_18 3.5355339059327378
E_p_18 nts_p_18 0 p18 0 0.07071067811865475
E_n_18 0 nt_n_18 nt_p_18 0 1
* Current sensor on center node for transfer to port 18
V_c_18 nt_c_18 0 0
* Transfer network from port 1 to port 18
R18_1 nt_n_1 nt_c_18 0.003124999999999963
X1837 nt_n_1 nt_c_18 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1838 nt_p_1 nt_c_18 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1839 nt_p_1 nt_c_18 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1840 nt_p_1 nt_c_18 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1841 nt_n_1 nt_c_18 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1842 nt_n_1 nt_c_18 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 2 to port 18
R18_2 nt_n_2 nt_c_18 0.003124999999999963
X1843 nt_n_2 nt_c_18 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1844 nt_p_2 nt_c_18 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1845 nt_p_2 nt_c_18 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1846 nt_p_2 nt_c_18 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1847 nt_n_2 nt_c_18 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1848 nt_n_2 nt_c_18 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 3 to port 18
R18_3 nt_n_3 nt_c_18 0.003124999999999963
X1849 nt_n_3 nt_c_18 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1850 nt_p_3 nt_c_18 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1851 nt_p_3 nt_c_18 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1852 nt_p_3 nt_c_18 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1853 nt_n_3 nt_c_18 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1854 nt_n_3 nt_c_18 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 4 to port 18
R18_4 nt_n_4 nt_c_18 0.003124999999999963
X1855 nt_n_4 nt_c_18 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1856 nt_p_4 nt_c_18 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1857 nt_p_4 nt_c_18 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1858 nt_p_4 nt_c_18 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1859 nt_n_4 nt_c_18 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1860 nt_n_4 nt_c_18 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 5 to port 18
R18_5 nt_n_5 nt_c_18 0.003124999999999963
X1861 nt_n_5 nt_c_18 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1862 nt_p_5 nt_c_18 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1863 nt_p_5 nt_c_18 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1864 nt_p_5 nt_c_18 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1865 nt_n_5 nt_c_18 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1866 nt_n_5 nt_c_18 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 6 to port 18
R18_6 nt_n_6 nt_c_18 0.003124999999999963
X1867 nt_n_6 nt_c_18 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1868 nt_p_6 nt_c_18 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1869 nt_p_6 nt_c_18 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1870 nt_p_6 nt_c_18 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1871 nt_n_6 nt_c_18 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1872 nt_n_6 nt_c_18 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 7 to port 18
R18_7 nt_n_7 nt_c_18 0.003124999999999963
X1873 nt_n_7 nt_c_18 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1874 nt_p_7 nt_c_18 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1875 nt_p_7 nt_c_18 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1876 nt_p_7 nt_c_18 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1877 nt_n_7 nt_c_18 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1878 nt_n_7 nt_c_18 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 8 to port 18
R18_8 nt_n_8 nt_c_18 0.003124999999999963
X1879 nt_n_8 nt_c_18 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1880 nt_p_8 nt_c_18 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1881 nt_p_8 nt_c_18 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1882 nt_p_8 nt_c_18 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1883 nt_n_8 nt_c_18 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1884 nt_n_8 nt_c_18 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 9 to port 18
R18_9 nt_n_9 nt_c_18 0.003124999999999963
X1885 nt_n_9 nt_c_18 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1886 nt_p_9 nt_c_18 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1887 nt_p_9 nt_c_18 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1888 nt_p_9 nt_c_18 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1889 nt_n_9 nt_c_18 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1890 nt_n_9 nt_c_18 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 10 to port 18
R18_10 nt_n_10 nt_c_18 0.003124999999999963
X1891 nt_n_10 nt_c_18 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1892 nt_p_10 nt_c_18 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1893 nt_p_10 nt_c_18 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1894 nt_p_10 nt_c_18 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1895 nt_n_10 nt_c_18 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1896 nt_n_10 nt_c_18 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 11 to port 18
R18_11 nt_n_11 nt_c_18 0.003124999999999963
X1897 nt_n_11 nt_c_18 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1898 nt_p_11 nt_c_18 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1899 nt_p_11 nt_c_18 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1900 nt_p_11 nt_c_18 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1901 nt_n_11 nt_c_18 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1902 nt_n_11 nt_c_18 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 12 to port 18
R18_12 nt_n_12 nt_c_18 0.003124999999999963
X1903 nt_n_12 nt_c_18 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1904 nt_p_12 nt_c_18 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1905 nt_p_12 nt_c_18 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1906 nt_p_12 nt_c_18 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1907 nt_n_12 nt_c_18 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1908 nt_n_12 nt_c_18 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 13 to port 18
R18_13 nt_n_13 nt_c_18 0.003124999999999963
X1909 nt_n_13 nt_c_18 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1910 nt_p_13 nt_c_18 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1911 nt_p_13 nt_c_18 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1912 nt_p_13 nt_c_18 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1913 nt_n_13 nt_c_18 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1914 nt_n_13 nt_c_18 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 14 to port 18
R18_14 nt_n_14 nt_c_18 0.003124999999999963
X1915 nt_n_14 nt_c_18 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1916 nt_p_14 nt_c_18 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1917 nt_p_14 nt_c_18 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1918 nt_p_14 nt_c_18 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1919 nt_n_14 nt_c_18 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1920 nt_n_14 nt_c_18 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 15 to port 18
R18_15 nt_n_15 nt_c_18 0.003124999999999963
X1921 nt_n_15 nt_c_18 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1922 nt_p_15 nt_c_18 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1923 nt_p_15 nt_c_18 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1924 nt_p_15 nt_c_18 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1925 nt_n_15 nt_c_18 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1926 nt_n_15 nt_c_18 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 16 to port 18
R18_16 nt_n_16 nt_c_18 0.003124999999999963
X1927 nt_n_16 nt_c_18 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1928 nt_p_16 nt_c_18 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1929 nt_p_16 nt_c_18 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1930 nt_p_16 nt_c_18 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1931 nt_n_16 nt_c_18 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1932 nt_n_16 nt_c_18 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 17 to port 18
R18_17 nt_n_17 nt_c_18 0.003124999999999963
X1933 nt_n_17 nt_c_18 rl_admittance res=2.7733601307884586e+17 ind=0.05119886123842035
X1934 nt_p_17 nt_c_18 rl_admittance res=187800143092.54297 ind=8.409869753766284
X1935 nt_p_17 nt_c_18 rl_admittance res=2830864960247.9546 ind=400.6893238451989
X1936 nt_p_17 nt_c_18 rl_admittance res=63732557064.23586 ind=35.261662271871394
X1937 nt_n_17 nt_c_18 rl_admittance res=112799484372.98152 ind=31.919389834390056
X1938 nt_n_17 nt_c_18 rl_admittance res=51262611157.92125 ind=93.72728905498322
* Transfer network from port 18 to port 18
R18_18 nt_p_18 nt_c_18 0.0007564900050830436
X1939 nt_p_18 nt_c_18 rl_admittance res=6.713812060922877e+16 ind=0.01239433452121846
X1940 nt_n_18 nt_c_18 rl_admittance res=0.00045787217518182793 ind=2.0503953265122565e-14
X1941 nt_p_18 nt_c_18 rl_admittance res=0.00054254751817662 ind=7.679384261163742e-14
X1942 nt_p_18 nt_c_18 rl_admittance res=0.0005564228350387422 ind=3.0785512135842906e-13
X1943 nt_n_18 nt_c_18 rl_admittance res=0.0005055304090704312 ind=1.4305226916553906e-13
X1944 nt_n_18 nt_c_18 rl_admittance res=0.00047272890640632993 ind=8.643258284073119e-13
.ENDS s_equivalent

.SUBCKT rcl_vccs_admittance n_pos n_neg res=1e3 cap=1e-9 ind=100e-12 gm=1e-3
L1 n_pos 1 {ind}
C1 1 2 {cap}
R1 2 n_neg {res}
G1 n_pos n_neg 1 2 {gm}
.ENDS rcl_vccs_admittance

.SUBCKT rl_admittance n_pos n_neg res=1e3 ind=100e-12
L1 n_pos 1 {ind}
R1 1 n_neg {res}
.ENDS rl_admittance

