* EQUIVALENT CIRCUIT FOR VECTOR FITTED
* Created by wyz
*
.SUBCKT s_equivalent p1 p2
*
* Port network for port 1
V1 p1 s1 0
R1 s1 0 50.0
Gd1_1 0 s1 p1 0 -0.019051175665602813
Fd1_1 0 s1 V1 -0.9525587832801408
Gr1_1_1 0 s1 x1_a1 0 22218617122.836678
Gr2_re_1_1 0 s1 x2_re_a1 0 34980203132.210045
Gr2_im_1_1 0 s1 x2_im_a1 0 52870233832.79671
Gr3_re_1_1 0 s1 x3_re_a1 0 69550148.1324326
Gr3_im_1_1 0 s1 x3_im_a1 0 -295109001.2402495
Gr4_re_1_1 0 s1 x4_re_a1 0 -132642686.58072104
Gr4_im_1_1 0 s1 x4_im_a1 0 -187312273.92280382
Gr5_re_1_1 0 s1 x5_re_a1 0 -91644162.8995502
Gr5_im_1_1 0 s1 x5_im_a1 0 -481749825.24265957
Gd1_2 0 s1 p2 0 3.9993436022022085e-05
Fd1_2 0 s1 V2 0.0019996718011011045
Gr1_1_2 0 s1 x1_a2 0 -16193390.35189798
Gr2_re_1_2 0 s1 x2_re_a2 0 -45811441.278188124
Gr2_im_1_2 0 s1 x2_im_a2 0 -9165465.085839208
Gr3_re_1_2 0 s1 x3_re_a2 0 60361226.284735784
Gr3_im_1_2 0 s1 x3_im_a2 0 -287683728.56018215
Gr4_re_1_2 0 s1 x4_re_a2 0 -138394278.02620646
Gr4_im_1_2 0 s1 x4_im_a2 0 -193103797.06061518
Gr5_re_1_2 0 s1 x5_re_a2 0 73029674.91777767
Gr5_im_1_2 0 s1 x5_im_a2 0 475538981.0820556
*
* State networks driven by port 1
Cx1_a1 x1_a1 0 1.0
Gx1_a1 0 x1_a1 p1 0 0.07071067811865475
Fx1_a1 0 x1_a1 V1 3.5355339059327378
Rp1_a1 0 x1_a1 4.027942112050941e-11
Cx2_re_a1 x2_re_a1 0 1.0
Gx2_re_a1 0 x2_re_a1 p1 0 0.1414213562373095
Fx2_re_a1 0 x2_re_a1 V1 7.0710678118654755
Rp2_re_re_a1 0 x2_re_a1 1.431065304142738e-11
Gp2_re_im_a1 0 x2_re_a1 x2_im_a1 0 97527973580.15533
Cx2_im_a1 x2_im_a1 0 1.0
Gp2_im_re_a1 0 x2_im_a1 x2_re_a1 0 -97527973580.15533
Rp2_im_im_a1 0 x2_im_a1 1.431065304142738e-11
Cx3_re_a1 x3_re_a1 0 1.0
Gx3_re_a1 0 x3_re_a1 p1 0 0.1414213562373095
Fx3_re_a1 0 x3_re_a1 V1 7.0710678118654755
Rp3_re_re_a1 0 x3_re_a1 1.099596071746407e-09
Gp3_re_im_a1 0 x3_re_a1 x3_im_a1 0 93663081207.82571
Cx3_im_a1 x3_im_a1 0 1.0
Gp3_im_re_a1 0 x3_im_a1 x3_re_a1 0 -93663081207.82571
Rp3_im_im_a1 0 x3_im_a1 1.099596071746407e-09
Cx4_re_a1 x4_re_a1 0 1.0
Gx4_re_a1 0 x4_re_a1 p1 0 0.1414213562373095
Fx4_re_a1 0 x4_re_a1 V1 7.0710678118654755
Rp4_re_re_a1 0 x4_re_a1 1.3403412255684957e-09
Gp4_re_im_a1 0 x4_re_a1 x4_im_a1 0 90484232971.93242
Cx4_im_a1 x4_im_a1 0 1.0
Gp4_im_re_a1 0 x4_im_a1 x4_re_a1 0 -90484232971.93242
Rp4_im_im_a1 0 x4_im_a1 1.3403412255684957e-09
Cx5_re_a1 x5_re_a1 0 1.0
Gx5_re_a1 0 x5_re_a1 p1 0 0.1414213562373095
Fx5_re_a1 0 x5_re_a1 V1 7.0710678118654755
Rp5_re_re_a1 0 x5_re_a1 6.178299898394442e-10
Gp5_re_im_a1 0 x5_re_a1 x5_im_a1 0 91963690751.78857
Cx5_im_a1 x5_im_a1 0 1.0
Gp5_im_re_a1 0 x5_im_a1 x5_re_a1 0 -91963690751.78857
Rp5_im_im_a1 0 x5_im_a1 6.178299898394442e-10
*
* Port network for port 2
V2 p2 s2 0
R2 s2 0 50.0
Gd2_1 0 s2 p1 0 3.999343602209308e-05
Fd2_1 0 s2 V1 0.001999671801104654
Gr1_2_1 0 s2 x1_a1 0 -16193390.352031434
Gr2_re_2_1 0 s2 x2_re_a1 0 -45811441.27827804
Gr2_im_2_1 0 s2 x2_im_a1 0 -9165465.08597713
Gr3_re_2_1 0 s2 x3_re_a1 0 60361226.284735724
Gr3_im_2_1 0 s2 x3_im_a1 0 -287683728.56018233
Gr4_re_2_1 0 s2 x4_re_a1 0 -138394278.0262065
Gr4_im_2_1 0 s2 x4_im_a1 0 -193103797.06061524
Gr5_re_2_1 0 s2 x5_re_a1 0 73029674.91777773
Gr5_im_2_1 0 s2 x5_im_a1 0 475538981.08205676
Gd2_2 0 s2 p2 0 -0.018964680676940113
Fd2_2 0 s2 V2 -0.9482340338470057
Gr1_2_2 0 s2 x1_a2 0 22195810474.297077
Gr2_re_2_2 0 s2 x2_re_a2 0 34845629036.36019
Gr2_im_2_2 0 s2 x2_im_a2 0 52777754102.26072
Gr3_re_2_2 0 s2 x3_re_a2 0 51845974.33171394
Gr3_im_2_2 0 s2 x3_im_a2 0 -280218053.0370414
Gr4_re_2_2 0 s2 x4_re_a2 0 -144502788.06752324
Gr4_im_2_2 0 s2 x4_im_a2 0 -198813279.71363327
Gr5_re_2_2 0 s2 x5_re_a2 0 -56294579.28884109
Gr5_im_2_2 0 s2 x5_im_a2 0 -470760867.0625005
*
* State networks driven by port 2
Cx1_a2 x1_a2 0 1.0
Gx1_a2 0 x1_a2 p2 0 0.07071067811865475
Fx1_a2 0 x1_a2 V2 3.5355339059327378
Rp1_a2 0 x1_a2 4.027942112050941e-11
Cx2_re_a2 x2_re_a2 0 1.0
Gx2_re_a2 0 x2_re_a2 p2 0 0.1414213562373095
Fx2_re_a2 0 x2_re_a2 V2 7.0710678118654755
Rp2_re_re_a2 0 x2_re_a2 1.431065304142738e-11
Gp2_re_im_a2 0 x2_re_a2 x2_im_a2 0 97527973580.15533
Cx2_im_a2 x2_im_a2 0 1.0
Gp2_im_re_a2 0 x2_im_a2 x2_re_a2 0 -97527973580.15533
Rp2_im_im_a2 0 x2_im_a2 1.431065304142738e-11
Cx3_re_a2 x3_re_a2 0 1.0
Gx3_re_a2 0 x3_re_a2 p2 0 0.1414213562373095
Fx3_re_a2 0 x3_re_a2 V2 7.0710678118654755
Rp3_re_re_a2 0 x3_re_a2 1.099596071746407e-09
Gp3_re_im_a2 0 x3_re_a2 x3_im_a2 0 93663081207.82571
Cx3_im_a2 x3_im_a2 0 1.0
Gp3_im_re_a2 0 x3_im_a2 x3_re_a2 0 -93663081207.82571
Rp3_im_im_a2 0 x3_im_a2 1.099596071746407e-09
Cx4_re_a2 x4_re_a2 0 1.0
Gx4_re_a2 0 x4_re_a2 p2 0 0.1414213562373095
Fx4_re_a2 0 x4_re_a2 V2 7.0710678118654755
Rp4_re_re_a2 0 x4_re_a2 1.3403412255684957e-09
Gp4_re_im_a2 0 x4_re_a2 x4_im_a2 0 90484232971.93242
Cx4_im_a2 x4_im_a2 0 1.0
Gp4_im_re_a2 0 x4_im_a2 x4_re_a2 0 -90484232971.93242
Rp4_im_im_a2 0 x4_im_a2 1.3403412255684957e-09
Cx5_re_a2 x5_re_a2 0 1.0
Gx5_re_a2 0 x5_re_a2 p2 0 0.1414213562373095
Fx5_re_a2 0 x5_re_a2 V2 7.0710678118654755
Rp5_re_re_a2 0 x5_re_a2 6.178299898394442e-10
Gp5_re_im_a2 0 x5_re_a2 x5_im_a2 0 91963690751.78857
Cx5_im_a2 x5_im_a2 0 1.0
Gp5_im_re_a2 0 x5_im_a2 x5_re_a2 0 -91963690751.78857
Rp5_im_im_a2 0 x5_im_a2 6.178299898394442e-10
.ENDS s_equivalent
